# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai31_1 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 3.85 5.55 4.1 8.3 ;
        RECT 1.05 5.55 1.3 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 2.25 0 2.5 1.6 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.95 2.95 1.45 3.25 ;
      LAYER Metal2 ;
        RECT 0.95 2.9 1.45 3.3 ;
      LAYER Via1 ;
        RECT 1.07 2.97 1.33 3.23 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 2.95 2.3 3.25 ;
      LAYER Metal2 ;
        RECT 1.8 2.9 2.3 3.3 ;
      LAYER Via1 ;
        RECT 1.92 2.97 2.18 3.23 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.55 4.25 3.05 4.55 ;
      LAYER Metal2 ;
        RECT 2.55 4.2 3.05 4.6 ;
      LAYER Via1 ;
        RECT 2.67 4.27 2.93 4.53 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 2.95 3.6 3.25 ;
      LAYER Metal2 ;
        RECT 3.1 2.9 3.6 3.3 ;
      LAYER Via1 ;
        RECT 3.22 2.97 3.48 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 4.9 4.25 5.2 ;
        RECT 3.95 1.05 4.2 2.6 ;
        RECT 3.85 2.35 4.1 5.2 ;
        RECT 3 4.9 3.25 7.25 ;
      LAYER Metal2 ;
        RECT 3.75 4.85 4.25 5.25 ;
      LAYER Via1 ;
        RECT 3.87 4.92 4.13 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.85 3.35 2.1 ;
      RECT 3.1 1.05 3.35 2.1 ;
      RECT 1.4 1.05 1.65 2.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai31_1
