# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__or2_1 0 0 ;
  SIZE 3.8 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 3.8 6.35 ;
        RECT 1.95 4.4 2.35 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.8 0.7 ;
        RECT 2.1 0 2.35 1.9 ;
        RECT 0.4 0 0.65 1.55 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.9 2.3 1.4 2.6 ;
      LAYER Metal2 ;
        RECT 0.9 2.25 1.4 2.65 ;
      LAYER Via1 ;
        RECT 1.02 2.32 1.28 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.65 2.95 2.15 3.25 ;
      LAYER Metal2 ;
        RECT 1.65 2.9 2.15 3.3 ;
      LAYER Via1 ;
        RECT 1.77 2.97 2.03 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.95 1.55 3.45 1.85 ;
        RECT 2.95 1.05 3.2 1.9 ;
        RECT 2.95 3.6 3.45 3.9 ;
        RECT 2.95 3.6 3.2 5.3 ;
      LAYER Metal2 ;
        RECT 2.95 3.55 3.45 3.95 ;
        RECT 2.95 1.5 3.45 1.9 ;
        RECT 3.05 1.5 3.35 3.95 ;
      LAYER Via1 ;
        RECT 3.07 3.62 3.33 3.88 ;
        RECT 3.07 1.57 3.33 1.83 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 3.05 0.8 5.3 ;
      RECT 0.55 3.85 2.7 4.15 ;
      RECT 2.4 3.05 2.7 4.15 ;
      RECT 2.4 3.05 2.95 3.35 ;
      RECT 0.4 1.8 0.65 3.35 ;
      RECT 0.4 1.8 1.5 2.05 ;
      RECT 1.25 1.05 1.5 2.05 ;
  END
END gf180mcu_osu_sc_gp9t3v3__or2_1
