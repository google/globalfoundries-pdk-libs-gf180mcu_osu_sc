* HSPICE file created from gf180mcu_osu_sc_12T_tiehi.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_tiehi Y
X0 Y a_19_11 VDD VDD pmos_3p3 w=34 l=6
X1 a_19_11 a_19_11 GND GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
