* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__clkbuf_16 A Y
X0 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X2 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X3 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X4 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X5 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X6 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X7 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X8 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X9 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X10 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X11 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X12 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X13 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X14 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X15 VSS A a_9_19 VSS nmos_3p3 w=17 l=6
X16 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X17 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X18 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X19 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X20 VSS a_9_19 Y VSS nmos_3p3 w=17 l=6
X21 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X22 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X23 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X24 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X25 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X26 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X27 Y a_9_19 VSS VSS nmos_3p3 w=17 l=6
X28 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X29 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X30 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
X31 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X32 Y a_9_19 VDD VDD pmos_3p3 w=34 l=6
X33 VDD a_9_19 Y VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
