# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffsrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsrn_1 0 0 ;
  SIZE 20.45 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 20.45 8.1 ;
        RECT 18.8 5.45 19.05 8.1 ;
        RECT 15.5 6.7 15.75 8.1 ;
        RECT 13.9 5.45 14.15 8.1 ;
        RECT 11.3 6.2 11.55 8.1 ;
        RECT 8.5 5.45 8.75 8.1 ;
        RECT 5.45 5.45 5.7 8.1 ;
        RECT 3.85 6.2 4.1 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 20.45 0.6 ;
        RECT 18.8 0 19.05 1.8 ;
        RECT 17.05 0 17.3 1.8 ;
        RECT 14.8 0 15.05 1.8 ;
        RECT 13.9 0 14.15 1.8 ;
        RECT 11.3 0 11.55 1.8 ;
        RECT 8.5 0 8.75 1.4 ;
        RECT 5.45 0 5.7 1.8 ;
        RECT 4.55 0 4.8 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 13.65 2.85 14.15 3.15 ;
      LAYER MET2 ;
        RECT 13.65 2.8 14.15 3.2 ;
      LAYER VIA12 ;
        RECT 13.77 2.87 14.03 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.95 3.5 6.45 3.8 ;
      LAYER MET2 ;
        RECT 5.95 3.45 6.45 3.85 ;
      LAYER VIA12 ;
        RECT 6.07 3.52 6.33 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 19.65 4.8 20.15 5.15 ;
        RECT 19.65 4.75 20.1 5.15 ;
        RECT 19.65 0.95 19.9 7.15 ;
      LAYER MET2 ;
        RECT 19.65 4.8 20.15 5.1 ;
        RECT 19.7 4.75 20.1 5.15 ;
      LAYER VIA12 ;
        RECT 19.77 4.82 20.03 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 17.95 4.15 19.4 4.45 ;
        RECT 19.05 2.05 19.3 4.45 ;
        RECT 17.95 2.05 19.3 2.3 ;
        RECT 17.95 4.15 18.2 7.15 ;
        RECT 17.95 0.95 18.2 2.3 ;
      LAYER MET2 ;
        RECT 18.9 4.15 19.4 4.45 ;
        RECT 18.95 4.1 19.35 4.5 ;
      LAYER VIA12 ;
        RECT 19.02 4.17 19.28 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.7 4.15 16.2 4.45 ;
        RECT 3.4 4.15 3.9 4.45 ;
      LAYER MET2 ;
        RECT 15.7 4.1 16.2 4.5 ;
        RECT 3.5 5.45 16.1 5.75 ;
        RECT 15.8 4.1 16.1 5.75 ;
        RECT 3.4 4.1 3.9 4.5 ;
        RECT 3.5 4.1 3.8 5.75 ;
      LAYER VIA12 ;
        RECT 3.52 4.17 3.78 4.43 ;
        RECT 15.82 4.17 16.08 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 18.2 2.8 18.6 3.2 ;
      RECT 17.85 2.85 18.65 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 16.6 2.1 17.2 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 16.6 0.9 16.9 2.5 ;
      RECT 2.75 0.9 16.9 1.2 ;
      RECT 14.7 2.1 15.2 2.5 ;
      RECT 14.7 1.55 15.1 2.5 ;
      RECT 9.85 1.5 10.25 1.9 ;
      RECT 9.8 1.55 15.1 1.85 ;
      RECT 14.75 4.75 15.15 5.15 ;
      RECT 10.8 4.75 11.2 5.15 ;
      RECT 10.75 4.8 15.2 5.1 ;
      RECT 12.95 4.1 13.4 4.5 ;
      RECT 11.75 4.1 12.15 4.5 ;
      RECT 10.1 4.1 10.6 4.5 ;
      RECT 7.3 4.1 7.75 4.5 ;
      RECT 7.3 4.15 13.4 4.45 ;
      RECT 12.1 2.8 12.5 3.2 ;
      RECT 10.15 2.8 10.55 3.2 ;
      RECT 10.1 2.85 12.6 3.15 ;
      RECT 10.85 3.45 11.25 3.85 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 8.15 2.15 8.55 2.55 ;
      RECT 4.4 2.15 4.9 2.55 ;
      RECT 4.4 2.2 8.6 2.5 ;
      RECT 17.1 4.75 17.6 5.15 ;
      RECT 4.4 3.45 4.9 3.85 ;
    LAYER VIA12 ;
      RECT 18.27 2.87 18.53 3.13 ;
      RECT 17.22 4.82 17.48 5.08 ;
      RECT 16.82 2.17 17.08 2.43 ;
      RECT 14.82 2.17 15.08 2.43 ;
      RECT 14.82 4.82 15.08 5.08 ;
      RECT 13.02 4.17 13.28 4.43 ;
      RECT 12.17 2.87 12.43 3.13 ;
      RECT 11.82 4.17 12.08 4.43 ;
      RECT 10.92 3.52 11.18 3.78 ;
      RECT 10.87 4.82 11.13 5.08 ;
      RECT 10.22 2.87 10.48 3.13 ;
      RECT 10.22 4.17 10.48 4.43 ;
      RECT 9.92 1.57 10.18 1.83 ;
      RECT 8.22 2.22 8.48 2.48 ;
      RECT 7.42 4.17 7.68 4.43 ;
      RECT 4.52 2.22 4.78 2.48 ;
      RECT 4.52 3.52 4.78 3.78 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 17.2 2.85 17.45 7.15 ;
      RECT 14.8 4.7 15.1 5.2 ;
      RECT 14.8 4.8 17.6 5.1 ;
      RECT 16.2 2.85 18.65 3.15 ;
      RECT 16.2 0.95 16.45 3.15 ;
      RECT 16.35 6.2 16.6 7.15 ;
      RECT 14.65 6.2 14.9 7.15 ;
      RECT 14.65 6.2 16.6 6.45 ;
      RECT 13.05 0.95 13.3 7.15 ;
      RECT 13 1.7 13.3 5.55 ;
      RECT 12.95 4.15 13.4 4.45 ;
      RECT 12.15 4.75 12.4 7.15 ;
      RECT 12.15 4.75 12.7 5 ;
      RECT 12.45 3.55 12.7 5 ;
      RECT 12.15 2.75 12.45 3.8 ;
      RECT 12.15 0.95 12.4 3.8 ;
      RECT 10.75 4.8 11.25 5.1 ;
      RECT 10.85 3.5 11.15 5.1 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 9.55 4.15 10.6 4.45 ;
      RECT 9.55 2.15 9.85 4.45 ;
      RECT 9.45 2.15 9.95 2.45 ;
      RECT 9.9 5.95 10.15 7.15 ;
      RECT 9 5.95 10.15 6.2 ;
      RECT 9 3.45 9.25 6.2 ;
      RECT 8.95 1.6 9.2 3.7 ;
      RECT 8.95 1.6 10.3 1.85 ;
      RECT 9.9 1.55 10.3 1.85 ;
      RECT 9.9 0.95 10.15 1.85 ;
      RECT 8.1 4.8 8.6 5.1 ;
      RECT 8.2 2.2 8.5 5.1 ;
      RECT 8.1 2.2 8.6 2.5 ;
      RECT 6.65 4.15 7.8 4.45 ;
      RECT 7.4 2.2 7.7 4.45 ;
      RECT 7.3 2.2 7.8 2.5 ;
      RECT 7.1 4.95 7.35 7.15 ;
      RECT 5.45 4.95 7.35 5.2 ;
      RECT 5.45 2.25 5.7 5.2 ;
      RECT 4.4 3.5 5.7 3.8 ;
      RECT 5.45 2.25 6.45 2.5 ;
      RECT 6.05 1.55 6.45 2.5 ;
      RECT 6.05 1.55 7.35 1.8 ;
      RECT 7.1 0.95 7.35 1.8 ;
      RECT 4.7 5.7 4.95 7.15 ;
      RECT 3 5.7 3.25 7.15 ;
      RECT 3 5.7 4.95 5.95 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 4.5 2.15 4.75 2.55 ;
      RECT 3.15 2.2 4.9 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 16.7 2.15 17.2 2.45 ;
      RECT 14.7 2.15 15.2 2.45 ;
      RECT 11.7 4.15 12.2 4.45 ;
      RECT 10.1 2.85 10.6 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsrn_1
