magic
tech gf180mcuC
timestamp 1661875376
<< nwell >>
rect 0 61 56 123
<< nmos >>
rect 16 19 22 36
rect 33 19 39 36
<< pmos >>
rect 19 70 25 104
rect 30 70 36 104
<< ndiff >>
rect 6 34 16 36
rect 6 21 8 34
rect 13 21 16 34
rect 6 19 16 21
rect 22 34 33 36
rect 22 21 25 34
rect 30 21 33 34
rect 22 19 33 21
rect 39 34 49 36
rect 39 21 42 34
rect 47 21 49 34
rect 39 19 49 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 70 30 104
rect 36 102 46 104
rect 36 79 39 102
rect 44 79 46 102
rect 36 70 46 79
<< ndiffc >>
rect 8 21 13 34
rect 25 21 30 34
rect 42 21 47 34
<< pdiffc >>
rect 11 72 16 102
rect 39 79 44 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
<< polysilicon >>
rect 19 104 25 109
rect 30 104 36 109
rect 19 66 25 70
rect 16 61 25 66
rect 30 67 36 70
rect 30 65 39 67
rect 30 63 47 65
rect 30 61 39 63
rect 16 52 22 61
rect 8 50 22 52
rect 8 44 11 50
rect 17 44 22 50
rect 8 42 22 44
rect 16 36 22 42
rect 33 57 39 61
rect 45 57 47 63
rect 33 55 47 57
rect 33 36 39 55
rect 16 14 22 19
rect 33 14 39 19
<< polycontact >>
rect 11 44 17 50
rect 39 57 45 63
<< metal1 >>
rect 0 118 56 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 56 118
rect 0 111 56 112
rect 11 102 16 111
rect 39 102 44 104
rect 39 77 44 79
rect 25 76 44 77
rect 11 70 16 72
rect 23 70 25 76
rect 31 72 44 76
rect 31 70 33 72
rect 9 44 11 50
rect 17 44 19 50
rect 8 34 13 36
rect 8 12 13 21
rect 25 34 30 70
rect 37 57 39 63
rect 45 57 47 63
rect 25 19 30 21
rect 42 34 47 36
rect 42 12 47 21
rect 0 11 56 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 56 11
rect 0 0 56 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 25 70 31 76
rect 11 44 17 50
rect 39 57 45 63
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 10 111 18 112
rect 34 111 42 112
rect 23 76 33 77
rect 23 70 25 76
rect 31 70 33 76
rect 23 69 33 70
rect 37 63 47 64
rect 37 57 39 63
rect 45 57 47 63
rect 37 56 47 57
rect 9 50 19 51
rect 9 44 11 50
rect 17 44 19 50
rect 9 43 19 44
rect 10 11 18 12
rect 34 11 42 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 10 4 18 5
rect 34 4 42 5
<< labels >>
rlabel metal2 13 115 13 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 14 47 14 47 1 A
port 1 n
rlabel metal2 28 73 28 73 1 Y
port 2 n
rlabel metal2 42 60 42 60 1 B
port 3 n
<< end >>
