magic
tech gf180mcuC
timestamp 1660269772
<< nwell >>
rect -2 97 94 159
<< nmos >>
rect 17 16 23 33
rect 51 16 57 33
rect 68 16 74 33
<< pmos >>
rect 17 106 23 140
rect 51 106 57 140
rect 68 106 74 140
<< ndiff >>
rect 7 31 17 33
rect 7 18 9 31
rect 14 18 17 31
rect 7 16 17 18
rect 23 31 33 33
rect 23 18 26 31
rect 31 18 33 31
rect 23 16 33 18
rect 41 31 51 33
rect 41 18 43 31
rect 48 18 51 31
rect 41 16 51 18
rect 57 31 68 33
rect 57 18 60 31
rect 65 18 68 31
rect 57 16 68 18
rect 74 31 84 33
rect 74 18 77 31
rect 82 18 84 31
rect 74 16 84 18
<< pdiff >>
rect 7 138 17 140
rect 7 108 9 138
rect 14 108 17 138
rect 7 106 17 108
rect 23 138 33 140
rect 23 108 26 138
rect 31 108 33 138
rect 23 106 33 108
rect 41 138 51 140
rect 41 108 43 138
rect 48 108 51 138
rect 41 106 51 108
rect 57 138 68 140
rect 57 108 60 138
rect 65 108 68 138
rect 57 106 68 108
rect 74 138 84 140
rect 74 108 77 138
rect 82 108 84 138
rect 74 106 84 108
<< ndiffc >>
rect 9 18 14 31
rect 26 18 31 31
rect 43 18 48 31
rect 60 18 65 31
rect 77 18 82 31
<< pdiffc >>
rect 9 108 14 138
rect 26 108 31 138
rect 43 108 48 138
rect 60 108 65 138
rect 77 108 82 138
<< psubdiff >>
rect 7 7 17 9
rect 7 2 9 7
rect 14 2 17 7
rect 7 0 17 2
rect 31 7 41 9
rect 31 2 33 7
rect 38 2 41 7
rect 31 0 41 2
rect 55 7 65 9
rect 55 2 57 7
rect 62 2 65 7
rect 55 0 65 2
<< nsubdiff >>
rect 7 154 17 156
rect 7 149 9 154
rect 14 149 17 154
rect 7 147 17 149
rect 31 154 41 156
rect 31 149 33 154
rect 38 149 41 154
rect 31 147 41 149
rect 55 154 65 156
rect 55 149 57 154
rect 62 149 65 154
rect 55 147 65 149
<< psubdiffcont >>
rect 9 2 14 7
rect 33 2 38 7
rect 57 2 62 7
<< nsubdiffcont >>
rect 9 149 14 154
rect 33 149 38 154
rect 57 149 62 154
<< polysilicon >>
rect 17 140 23 145
rect 51 140 57 145
rect 68 140 74 145
rect 17 103 23 106
rect 51 103 57 106
rect 17 98 57 103
rect 17 62 23 98
rect 28 86 38 89
rect 68 86 74 106
rect 28 80 30 86
rect 36 80 74 86
rect 28 77 38 80
rect 10 60 23 62
rect 10 55 12 60
rect 17 55 74 60
rect 10 53 23 55
rect 17 33 23 53
rect 28 47 38 50
rect 28 41 30 47
rect 36 46 38 47
rect 36 41 57 46
rect 28 38 38 41
rect 51 33 57 41
rect 68 33 74 55
rect 17 11 23 16
rect 51 11 57 16
rect 68 11 74 16
<< polycontact >>
rect 30 80 36 86
rect 12 55 17 60
rect 30 41 36 47
<< metal1 >>
rect -2 154 94 159
rect -2 148 9 154
rect 15 148 33 154
rect 39 148 57 154
rect 63 148 94 154
rect -2 147 94 148
rect 9 138 14 147
rect 9 106 14 108
rect 26 138 31 140
rect 26 86 31 108
rect 43 138 48 140
rect 26 80 30 86
rect 36 80 38 86
rect 9 54 11 60
rect 17 54 19 60
rect 26 47 31 80
rect 43 74 48 108
rect 60 138 65 140
rect 60 100 65 108
rect 77 138 82 140
rect 58 99 68 100
rect 58 93 60 99
rect 66 93 68 99
rect 58 92 68 93
rect 43 73 55 74
rect 43 67 47 73
rect 53 67 55 73
rect 43 66 55 67
rect 26 41 30 47
rect 36 41 38 47
rect 9 31 14 33
rect 9 9 14 18
rect 26 31 31 41
rect 26 16 31 18
rect 43 31 48 66
rect 43 16 48 18
rect 60 31 65 92
rect 77 87 82 108
rect 73 86 83 87
rect 73 80 75 86
rect 81 80 83 86
rect 73 79 83 80
rect 60 16 65 18
rect 77 31 82 79
rect 77 16 82 18
rect -2 8 94 9
rect -2 2 9 8
rect 15 2 33 8
rect 39 2 57 8
rect 63 2 94 8
rect -2 -3 94 2
<< via1 >>
rect 9 149 14 154
rect 14 149 15 154
rect 9 148 15 149
rect 33 149 38 154
rect 38 149 39 154
rect 33 148 39 149
rect 57 149 62 154
rect 62 149 63 154
rect 57 148 63 149
rect 11 55 12 60
rect 12 55 17 60
rect 11 54 17 55
rect 60 93 66 99
rect 47 67 53 73
rect 75 80 81 86
rect 9 7 15 8
rect 9 2 14 7
rect 14 2 15 7
rect 33 7 39 8
rect 33 2 38 7
rect 38 2 39 7
rect 57 7 63 8
rect 57 2 62 7
rect 62 2 63 7
<< metal2 >>
rect 8 154 16 155
rect 32 154 40 155
rect 56 154 64 155
rect 7 148 9 154
rect 15 148 17 154
rect 31 148 33 154
rect 39 148 41 154
rect 55 148 57 154
rect 63 148 65 154
rect 8 147 16 148
rect 32 147 40 148
rect 56 147 64 148
rect 58 99 68 100
rect 58 93 60 99
rect 66 93 68 99
rect 58 92 68 93
rect 73 86 83 87
rect 73 80 75 86
rect 81 80 83 86
rect 73 79 83 80
rect 45 73 55 74
rect 45 67 47 73
rect 53 67 55 73
rect 45 66 55 67
rect 9 60 19 61
rect 9 54 11 60
rect 17 54 19 60
rect 9 53 19 54
rect 8 8 16 9
rect 32 8 40 9
rect 56 8 64 9
rect 7 2 9 8
rect 15 2 17 8
rect 31 2 33 8
rect 39 2 41 8
rect 55 2 57 8
rect 63 2 65 8
rect 8 1 16 2
rect 32 1 40 2
rect 56 1 64 2
<< labels >>
rlabel metal2 12 5 12 5 1 GND
rlabel metal2 12 151 12 151 1 VDD
rlabel metal2 63 96 63 96 1 Y
port 2 n
rlabel metal2 50 70 50 70 1 A
port 4 n
rlabel metal2 78 83 78 83 1 B
port 5 n
rlabel metal2 14 57 14 57 1 Sel
port 3 n
<< end >>
