magic
tech gf180mcuC
timestamp 1661874219
<< nwell >>
rect 0 61 290 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 57 19 63 36
rect 80 19 86 36
rect 91 19 97 36
rect 108 19 114 36
rect 119 19 125 36
rect 142 19 148 36
rect 163 19 169 36
rect 180 19 186 36
rect 216 19 222 36
rect 248 19 254 36
rect 265 19 271 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 57 70 63 104
rect 80 70 86 104
rect 91 70 97 104
rect 108 70 114 104
rect 119 70 125 104
rect 142 70 148 104
rect 163 70 169 104
rect 180 70 186 104
rect 216 70 222 104
rect 248 70 254 104
rect 265 70 271 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 27 36 36
rect 25 21 28 27
rect 33 21 36 27
rect 25 19 36 21
rect 42 19 57 36
rect 63 27 80 36
rect 63 21 66 27
rect 77 21 80 27
rect 63 19 80 21
rect 86 19 91 36
rect 97 26 108 36
rect 97 21 100 26
rect 105 21 108 26
rect 97 19 108 21
rect 114 19 119 36
rect 125 26 142 36
rect 125 21 128 26
rect 139 21 142 26
rect 125 19 142 21
rect 148 19 163 36
rect 169 27 180 36
rect 169 21 172 27
rect 177 21 180 27
rect 169 19 180 21
rect 186 26 196 36
rect 186 21 189 26
rect 194 21 196 26
rect 186 19 196 21
rect 206 26 216 36
rect 206 21 208 26
rect 213 21 216 26
rect 206 19 216 21
rect 222 34 232 36
rect 222 21 225 34
rect 230 21 232 34
rect 222 19 232 21
rect 238 34 248 36
rect 238 21 240 34
rect 245 21 248 34
rect 238 19 248 21
rect 254 30 265 36
rect 254 21 257 30
rect 262 21 265 30
rect 254 19 265 21
rect 271 34 281 36
rect 271 21 274 34
rect 279 21 281 34
rect 271 19 281 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 36 104
rect 25 97 28 102
rect 33 97 36 102
rect 25 70 36 97
rect 42 70 57 104
rect 63 102 80 104
rect 63 86 66 102
rect 77 86 80 102
rect 63 70 80 86
rect 86 70 91 104
rect 97 102 108 104
rect 97 84 100 102
rect 105 84 108 102
rect 97 70 108 84
rect 114 70 119 104
rect 125 102 142 104
rect 125 86 128 102
rect 139 86 142 102
rect 125 70 142 86
rect 148 70 163 104
rect 169 102 180 104
rect 169 97 172 102
rect 177 97 180 102
rect 169 70 180 97
rect 186 102 196 104
rect 186 72 189 102
rect 194 72 196 102
rect 186 70 196 72
rect 206 102 216 104
rect 206 72 208 102
rect 213 72 216 102
rect 206 70 216 72
rect 222 102 232 104
rect 222 72 225 102
rect 230 72 232 102
rect 222 70 232 72
rect 238 102 248 104
rect 238 72 240 102
rect 245 72 248 102
rect 238 70 248 72
rect 254 102 265 104
rect 254 83 257 102
rect 262 83 265 102
rect 254 70 265 83
rect 271 102 281 104
rect 271 89 274 102
rect 279 89 281 102
rect 271 70 281 89
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 27
rect 66 21 77 27
rect 100 21 105 26
rect 128 21 139 26
rect 172 21 177 27
rect 189 21 194 26
rect 208 21 213 26
rect 225 21 230 34
rect 240 21 245 34
rect 257 21 262 30
rect 274 21 279 34
<< pdiffc >>
rect 11 72 16 102
rect 28 97 33 102
rect 66 86 77 102
rect 100 84 105 102
rect 128 86 139 102
rect 172 97 177 102
rect 189 72 194 102
rect 208 72 213 102
rect 225 72 230 102
rect 240 72 245 102
rect 257 83 262 102
rect 274 89 279 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 129 10 138 12
rect 129 5 131 10
rect 136 5 138 10
rect 129 3 138 5
rect 153 10 162 12
rect 153 5 155 10
rect 160 5 162 10
rect 153 3 162 5
rect 177 10 186 12
rect 177 5 179 10
rect 184 5 186 10
rect 177 3 186 5
rect 201 10 210 12
rect 201 5 203 10
rect 208 5 210 10
rect 201 3 210 5
rect 225 10 234 12
rect 225 5 227 10
rect 232 5 234 10
rect 225 3 234 5
rect 249 10 258 12
rect 249 5 251 10
rect 256 5 258 10
rect 249 3 258 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
rect 81 118 90 120
rect 81 113 83 118
rect 88 113 90 118
rect 81 111 90 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
rect 129 118 138 120
rect 129 113 131 118
rect 136 113 138 118
rect 129 111 138 113
rect 153 118 162 120
rect 153 113 155 118
rect 160 113 162 118
rect 153 111 162 113
rect 177 118 186 120
rect 177 113 179 118
rect 184 113 186 118
rect 177 111 186 113
rect 201 118 210 120
rect 201 113 203 118
rect 208 113 210 118
rect 201 111 210 113
rect 225 118 234 120
rect 225 113 227 118
rect 232 113 234 118
rect 225 111 234 113
rect 249 118 258 120
rect 249 113 251 118
rect 256 113 258 118
rect 249 111 258 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
rect 131 5 136 10
rect 155 5 160 10
rect 179 5 184 10
rect 203 5 208 10
rect 227 5 232 10
rect 251 5 256 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
rect 107 113 112 118
rect 131 113 136 118
rect 155 113 160 118
rect 179 113 184 118
rect 203 113 208 118
rect 227 113 232 118
rect 251 113 256 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 57 104 63 109
rect 80 104 86 109
rect 91 104 97 109
rect 108 104 114 109
rect 119 104 125 109
rect 142 104 148 109
rect 163 104 169 109
rect 180 104 186 109
rect 216 104 222 109
rect 248 104 254 109
rect 265 104 271 109
rect 19 68 25 70
rect 19 66 29 68
rect 19 60 21 66
rect 27 60 29 66
rect 36 65 42 70
rect 57 68 63 70
rect 50 66 63 68
rect 19 58 29 60
rect 34 63 45 65
rect 19 36 25 58
rect 34 57 37 63
rect 43 57 45 63
rect 50 61 53 66
rect 58 65 63 66
rect 58 61 60 65
rect 50 59 60 61
rect 80 57 86 70
rect 91 68 97 70
rect 108 68 114 70
rect 91 61 114 68
rect 34 55 45 57
rect 36 36 42 55
rect 65 52 86 57
rect 65 48 71 52
rect 53 46 71 48
rect 99 47 105 61
rect 119 57 125 70
rect 142 68 148 70
rect 142 66 154 68
rect 142 65 146 66
rect 144 60 146 65
rect 152 60 154 66
rect 144 58 154 60
rect 119 52 139 57
rect 163 52 169 70
rect 180 65 186 70
rect 180 63 190 65
rect 180 57 182 63
rect 188 57 190 63
rect 216 59 222 70
rect 248 59 254 70
rect 180 55 190 57
rect 210 57 222 59
rect 134 50 139 52
rect 161 50 171 52
rect 53 40 56 46
rect 62 40 71 46
rect 76 45 86 47
rect 76 40 78 45
rect 84 40 86 45
rect 53 38 65 40
rect 76 38 86 40
rect 57 36 63 38
rect 80 36 86 38
rect 91 46 105 47
rect 91 45 114 46
rect 91 40 94 45
rect 100 40 114 45
rect 91 38 114 40
rect 91 36 97 38
rect 108 36 114 38
rect 119 45 129 47
rect 119 40 121 45
rect 127 40 129 45
rect 134 46 148 50
rect 134 40 139 46
rect 145 40 148 46
rect 161 44 163 50
rect 169 44 171 50
rect 161 42 171 44
rect 119 38 129 40
rect 137 38 148 40
rect 119 36 125 38
rect 142 36 148 38
rect 163 36 169 42
rect 180 36 186 55
rect 210 51 212 57
rect 218 51 222 57
rect 210 49 222 51
rect 243 57 254 59
rect 243 51 245 57
rect 251 51 254 57
rect 265 52 271 70
rect 243 49 254 51
rect 216 36 222 49
rect 248 36 254 49
rect 259 50 271 52
rect 259 44 261 50
rect 267 44 271 50
rect 259 42 271 44
rect 265 36 271 42
rect 19 14 25 19
rect 36 14 42 19
rect 57 14 63 19
rect 80 14 86 19
rect 91 14 97 19
rect 108 14 114 19
rect 119 14 125 19
rect 142 14 148 19
rect 163 14 169 19
rect 180 14 186 19
rect 216 14 222 19
rect 248 14 254 19
rect 265 14 271 19
<< polycontact >>
rect 21 60 27 66
rect 37 57 43 63
rect 53 61 58 66
rect 146 60 152 66
rect 182 57 188 63
rect 56 40 62 46
rect 78 40 84 45
rect 94 40 100 45
rect 121 40 127 45
rect 139 40 145 46
rect 163 44 169 50
rect 212 51 218 57
rect 245 51 251 57
rect 261 44 267 50
<< metal1 >>
rect 0 118 290 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 131 118
rect 137 112 155 118
rect 161 112 179 118
rect 185 112 203 118
rect 209 112 227 118
rect 233 112 251 118
rect 257 112 290 118
rect 0 111 290 112
rect 11 102 16 104
rect 28 102 33 111
rect 28 95 33 97
rect 66 102 77 104
rect 11 47 16 72
rect 10 46 16 47
rect 8 40 10 46
rect 10 38 16 40
rect 11 34 16 38
rect 21 86 66 90
rect 21 84 77 86
rect 100 102 105 111
rect 21 66 27 84
rect 100 82 105 84
rect 128 102 139 104
rect 172 102 177 111
rect 172 95 177 97
rect 189 102 194 104
rect 134 84 139 86
rect 161 84 163 90
rect 169 84 171 90
rect 128 82 134 84
rect 163 82 169 84
rect 208 102 213 111
rect 194 72 200 75
rect 189 70 200 72
rect 208 70 213 72
rect 225 102 230 104
rect 27 60 29 66
rect 21 41 27 60
rect 35 57 37 63
rect 43 57 45 63
rect 50 61 53 66
rect 58 61 146 66
rect 50 60 146 61
rect 152 65 179 66
rect 152 63 188 65
rect 152 60 182 63
rect 78 46 84 60
rect 94 46 100 47
rect 21 36 45 41
rect 54 40 56 46
rect 62 40 64 46
rect 76 45 86 46
rect 76 40 78 45
rect 84 40 86 45
rect 92 40 94 46
rect 100 40 102 46
rect 121 45 127 60
rect 180 57 182 60
rect 188 57 190 63
rect 195 50 200 70
rect 139 46 145 48
rect 119 40 121 45
rect 127 40 129 45
rect 138 40 139 46
rect 145 40 151 46
rect 161 44 163 50
rect 169 44 171 50
rect 189 44 200 50
rect 212 57 218 59
rect 119 39 129 40
rect 139 38 151 40
rect 40 33 45 36
rect 145 37 151 38
rect 11 19 16 21
rect 28 27 33 30
rect 40 28 77 33
rect 126 28 128 33
rect 28 12 33 21
rect 66 27 77 28
rect 66 19 77 21
rect 100 26 105 28
rect 100 12 105 21
rect 134 27 139 33
rect 145 29 151 31
rect 189 37 195 44
rect 212 39 218 51
rect 225 57 230 72
rect 240 102 245 104
rect 257 102 262 111
rect 257 81 262 83
rect 274 102 279 104
rect 279 89 285 90
rect 274 83 277 89
rect 283 83 285 89
rect 274 82 284 83
rect 245 72 261 76
rect 240 70 261 72
rect 267 70 269 76
rect 225 51 245 57
rect 251 51 253 57
rect 210 33 212 39
rect 218 33 220 39
rect 225 34 230 51
rect 261 50 267 70
rect 261 42 267 44
rect 128 26 139 27
rect 128 19 139 21
rect 172 27 177 30
rect 172 12 177 21
rect 189 29 195 31
rect 189 26 194 29
rect 189 19 194 21
rect 208 26 213 28
rect 208 12 213 21
rect 225 19 230 21
rect 240 37 267 42
rect 240 34 245 37
rect 274 34 279 82
rect 240 19 245 21
rect 257 30 262 32
rect 257 12 262 21
rect 274 19 279 21
rect 0 11 290 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 131 11
rect 137 5 155 11
rect 161 5 179 11
rect 185 5 203 11
rect 209 5 227 11
rect 233 5 251 11
rect 257 5 290 11
rect 0 0 290 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 131 113 136 118
rect 136 113 137 118
rect 131 112 137 113
rect 155 113 160 118
rect 160 113 161 118
rect 155 112 161 113
rect 179 113 184 118
rect 184 113 185 118
rect 179 112 185 113
rect 203 113 208 118
rect 208 113 209 118
rect 203 112 209 113
rect 227 113 232 118
rect 232 113 233 118
rect 227 112 233 113
rect 251 113 256 118
rect 256 113 257 118
rect 251 112 257 113
rect 10 40 16 46
rect 128 86 134 90
rect 128 84 134 86
rect 163 84 169 90
rect 37 57 43 63
rect 56 40 62 46
rect 94 45 100 46
rect 94 40 100 45
rect 182 57 188 63
rect 163 44 169 50
rect 128 27 134 33
rect 145 31 151 37
rect 277 83 283 89
rect 261 70 267 76
rect 245 51 251 57
rect 189 31 195 37
rect 212 33 218 39
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 131 10 137 11
rect 131 5 136 10
rect 136 5 137 10
rect 155 10 161 11
rect 155 5 160 10
rect 160 5 161 10
rect 179 10 185 11
rect 179 5 184 10
rect 184 5 185 10
rect 203 10 209 11
rect 203 5 208 10
rect 208 5 209 10
rect 227 10 233 11
rect 227 5 232 10
rect 232 5 233 10
rect 251 10 257 11
rect 251 5 256 10
rect 256 5 257 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 129 112 131 118
rect 137 112 139 118
rect 153 112 155 118
rect 161 112 163 118
rect 177 112 179 118
rect 185 112 187 118
rect 201 112 203 118
rect 209 112 211 118
rect 225 112 227 118
rect 233 112 235 118
rect 249 112 251 118
rect 257 112 259 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 56 98 151 104
rect 35 63 45 64
rect 34 57 37 63
rect 43 57 46 63
rect 35 56 45 57
rect 56 47 62 98
rect 128 91 134 92
rect 127 90 135 91
rect 127 84 128 90
rect 134 84 135 90
rect 127 83 135 84
rect 9 46 17 47
rect 55 46 64 47
rect 93 46 101 47
rect 8 40 10 46
rect 16 40 18 46
rect 54 40 56 46
rect 62 40 64 46
rect 92 40 94 46
rect 100 40 102 46
rect 9 39 17 40
rect 55 39 64 40
rect 93 39 101 40
rect 10 27 16 39
rect 94 27 100 39
rect 128 34 134 83
rect 145 38 151 98
rect 162 90 170 91
rect 161 84 163 90
rect 169 84 229 90
rect 276 89 284 90
rect 162 83 170 84
rect 163 51 169 83
rect 181 63 189 64
rect 180 57 182 63
rect 188 57 190 63
rect 223 57 229 84
rect 275 83 277 89
rect 283 83 285 89
rect 276 82 284 83
rect 260 76 268 77
rect 259 70 261 76
rect 267 70 269 76
rect 260 69 268 70
rect 244 57 252 58
rect 181 56 189 57
rect 223 51 245 57
rect 251 51 253 57
rect 162 50 170 51
rect 244 50 252 51
rect 161 44 163 50
rect 169 44 171 50
rect 162 43 170 44
rect 211 39 219 40
rect 144 37 152 38
rect 188 37 196 38
rect 127 33 135 34
rect 126 27 128 33
rect 134 27 135 33
rect 143 31 145 37
rect 151 31 189 37
rect 195 31 198 37
rect 204 33 212 39
rect 218 33 220 39
rect 204 32 219 33
rect 144 30 152 31
rect 188 30 196 31
rect 10 21 100 27
rect 127 26 135 27
rect 128 24 135 26
rect 204 24 210 32
rect 128 18 210 24
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 129 5 131 11
rect 137 5 139 11
rect 153 5 155 11
rect 161 5 163 11
rect 177 5 179 11
rect 185 5 187 11
rect 201 5 203 11
rect 209 5 211 11
rect 225 5 227 11
rect 233 5 235 11
rect 249 5 251 11
rect 257 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 13 8 13 8 1 GND
rlabel metal2 40 60 40 60 1 D
port 1 n
rlabel metal2 185 60 185 60 1 CLK
port 6 n
rlabel metal2 280 86 280 86 1 Q
port 4 n
rlabel metal2 264 73 264 73 1 QN
port 5 n
<< end >>
