magic
tech gf180mcuC
timestamp 1661888053
<< nwell >>
rect 0 61 410 123
<< nmos >>
rect 19 19 25 36
rect 54 19 60 36
rect 71 19 77 36
rect 82 19 88 36
rect 122 19 128 36
rect 143 19 149 36
rect 166 19 172 36
rect 177 19 183 36
rect 194 19 200 36
rect 205 19 211 36
rect 228 19 234 36
rect 249 19 255 36
rect 266 19 272 36
rect 304 19 310 36
rect 315 19 321 36
rect 332 19 338 36
rect 367 19 373 36
rect 384 19 390 36
<< pmos >>
rect 19 70 25 104
rect 51 70 57 104
rect 68 70 74 104
rect 85 70 91 104
rect 122 70 128 104
rect 143 70 149 104
rect 166 70 172 104
rect 177 70 183 104
rect 194 70 200 104
rect 205 70 211 104
rect 228 70 234 104
rect 249 70 255 104
rect 266 70 272 104
rect 301 70 307 104
rect 318 70 324 104
rect 335 70 341 104
rect 367 70 373 104
rect 384 70 390 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 35 36
rect 25 21 28 34
rect 33 21 35 34
rect 25 19 35 21
rect 44 26 54 36
rect 44 21 46 26
rect 51 21 54 26
rect 44 19 54 21
rect 60 31 71 36
rect 60 21 63 31
rect 68 21 71 31
rect 60 19 71 21
rect 77 19 82 36
rect 88 27 98 36
rect 88 21 91 27
rect 96 21 98 27
rect 88 19 98 21
rect 112 27 122 36
rect 112 21 114 27
rect 119 21 122 27
rect 112 19 122 21
rect 128 19 143 36
rect 149 27 166 36
rect 149 21 152 27
rect 163 21 166 27
rect 149 19 166 21
rect 172 19 177 36
rect 183 26 194 36
rect 183 21 186 26
rect 191 21 194 26
rect 183 19 194 21
rect 200 19 205 36
rect 211 26 228 36
rect 211 21 214 26
rect 225 21 228 26
rect 211 19 228 21
rect 234 19 249 36
rect 255 31 266 36
rect 255 21 258 31
rect 263 21 266 31
rect 255 19 266 21
rect 272 34 282 36
rect 272 21 275 34
rect 280 21 282 34
rect 272 19 282 21
rect 294 34 304 36
rect 294 21 296 34
rect 301 21 304 34
rect 294 19 304 21
rect 310 19 315 36
rect 321 29 332 36
rect 321 21 324 29
rect 329 21 332 29
rect 321 19 332 21
rect 338 26 348 36
rect 338 21 341 26
rect 346 21 348 26
rect 338 19 348 21
rect 357 34 367 36
rect 357 21 359 34
rect 364 21 367 34
rect 357 19 367 21
rect 373 30 384 36
rect 373 21 376 30
rect 381 21 384 30
rect 373 19 384 21
rect 390 34 400 36
rect 390 21 393 34
rect 398 21 400 34
rect 390 19 400 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 35 104
rect 25 72 28 102
rect 33 72 35 102
rect 25 70 35 72
rect 41 102 51 104
rect 41 88 43 102
rect 48 88 51 102
rect 41 70 51 88
rect 57 102 68 104
rect 57 87 60 102
rect 65 87 68 102
rect 57 70 68 87
rect 74 102 85 104
rect 74 87 77 102
rect 82 87 85 102
rect 74 70 85 87
rect 91 102 101 104
rect 91 87 94 102
rect 99 87 101 102
rect 91 70 101 87
rect 112 102 122 104
rect 112 97 114 102
rect 119 97 122 102
rect 112 70 122 97
rect 128 70 143 104
rect 149 102 166 104
rect 149 86 152 102
rect 163 86 166 102
rect 149 70 166 86
rect 172 70 177 104
rect 183 102 194 104
rect 183 84 186 102
rect 191 84 194 102
rect 183 70 194 84
rect 200 70 205 104
rect 211 102 228 104
rect 211 76 214 102
rect 225 76 228 102
rect 211 70 228 76
rect 234 70 249 104
rect 255 102 266 104
rect 255 97 258 102
rect 263 97 266 102
rect 255 70 266 97
rect 272 102 282 104
rect 272 74 275 102
rect 280 74 282 102
rect 272 70 282 74
rect 291 102 301 104
rect 291 87 293 102
rect 298 87 301 102
rect 291 70 301 87
rect 307 102 318 104
rect 307 87 310 102
rect 315 87 318 102
rect 307 70 318 87
rect 324 102 335 104
rect 324 87 327 102
rect 332 87 335 102
rect 324 70 335 87
rect 341 102 351 104
rect 341 88 344 102
rect 349 88 351 102
rect 341 70 351 88
rect 357 102 367 104
rect 357 73 359 102
rect 364 73 367 102
rect 357 70 367 73
rect 373 102 384 104
rect 373 83 376 102
rect 381 83 384 102
rect 373 70 384 83
rect 390 102 400 104
rect 390 72 393 102
rect 398 72 400 102
rect 390 70 400 72
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 46 21 51 26
rect 63 21 68 31
rect 91 21 96 27
rect 114 21 119 27
rect 152 21 163 27
rect 186 21 191 26
rect 214 21 225 26
rect 258 21 263 31
rect 275 21 280 34
rect 296 21 301 34
rect 324 21 329 29
rect 341 21 346 26
rect 359 21 364 34
rect 376 21 381 30
rect 393 21 398 34
<< pdiffc >>
rect 11 72 16 102
rect 28 72 33 102
rect 43 88 48 102
rect 60 87 65 102
rect 77 87 82 102
rect 94 87 99 102
rect 114 97 119 102
rect 152 86 163 102
rect 186 84 191 102
rect 214 76 225 102
rect 258 97 263 102
rect 275 74 280 102
rect 293 87 298 102
rect 310 87 315 102
rect 327 87 332 102
rect 344 88 349 102
rect 359 73 364 102
rect 376 83 381 102
rect 393 72 398 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 34 10 43 12
rect 34 5 36 10
rect 41 5 43 10
rect 34 3 43 5
rect 58 10 67 12
rect 58 5 60 10
rect 65 5 67 10
rect 58 3 67 5
rect 82 10 91 12
rect 82 5 84 10
rect 89 5 91 10
rect 82 3 91 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 129 10 138 12
rect 129 5 131 10
rect 136 5 138 10
rect 129 3 138 5
rect 153 10 162 12
rect 153 5 155 10
rect 160 5 162 10
rect 153 3 162 5
rect 177 10 186 12
rect 177 5 179 10
rect 184 5 186 10
rect 177 3 186 5
rect 201 10 210 12
rect 201 5 203 10
rect 208 5 210 10
rect 201 3 210 5
rect 225 10 234 12
rect 225 5 227 10
rect 232 5 234 10
rect 225 3 234 5
rect 249 10 258 12
rect 249 5 251 10
rect 256 5 258 10
rect 249 3 258 5
rect 273 10 282 12
rect 273 5 275 10
rect 280 5 282 10
rect 273 3 282 5
rect 297 10 306 12
rect 297 5 299 10
rect 304 5 306 10
rect 297 3 306 5
rect 321 10 330 12
rect 321 5 323 10
rect 328 5 330 10
rect 321 3 330 5
rect 345 10 354 12
rect 345 5 347 10
rect 352 5 354 10
rect 345 3 354 5
rect 369 10 378 12
rect 369 5 371 10
rect 376 5 378 10
rect 369 3 378 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 34 118 43 120
rect 34 113 36 118
rect 41 113 43 118
rect 34 111 43 113
rect 58 118 67 120
rect 58 113 60 118
rect 65 113 67 118
rect 58 111 67 113
rect 82 118 91 120
rect 82 113 84 118
rect 89 113 91 118
rect 82 111 91 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
rect 129 118 138 120
rect 129 113 131 118
rect 136 113 138 118
rect 129 111 138 113
rect 153 118 162 120
rect 153 113 155 118
rect 160 113 162 118
rect 153 111 162 113
rect 177 118 186 120
rect 177 113 179 118
rect 184 113 186 118
rect 177 111 186 113
rect 201 118 210 120
rect 201 113 203 118
rect 208 113 210 118
rect 201 111 210 113
rect 225 118 234 120
rect 225 113 227 118
rect 232 113 234 118
rect 225 111 234 113
rect 249 118 258 120
rect 249 113 251 118
rect 256 113 258 118
rect 249 111 258 113
rect 273 118 282 120
rect 273 113 275 118
rect 280 113 282 118
rect 273 111 282 113
rect 297 118 306 120
rect 297 113 299 118
rect 304 113 306 118
rect 297 111 306 113
rect 321 118 330 120
rect 321 113 323 118
rect 328 113 330 118
rect 321 111 330 113
rect 345 118 354 120
rect 345 113 347 118
rect 352 113 354 118
rect 345 111 354 113
rect 369 118 378 120
rect 369 113 371 118
rect 376 113 378 118
rect 369 111 378 113
<< psubdiffcont >>
rect 11 5 16 10
rect 36 5 41 10
rect 60 5 65 10
rect 84 5 89 10
rect 107 5 112 10
rect 131 5 136 10
rect 155 5 160 10
rect 179 5 184 10
rect 203 5 208 10
rect 227 5 232 10
rect 251 5 256 10
rect 275 5 280 10
rect 299 5 304 10
rect 323 5 328 10
rect 347 5 352 10
rect 371 5 376 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 36 113 41 118
rect 60 113 65 118
rect 84 113 89 118
rect 107 113 112 118
rect 131 113 136 118
rect 155 113 160 118
rect 179 113 184 118
rect 203 113 208 118
rect 227 113 232 118
rect 251 113 256 118
rect 275 113 280 118
rect 299 113 304 118
rect 323 113 328 118
rect 347 113 352 118
rect 371 113 376 118
<< polysilicon >>
rect 19 104 25 109
rect 51 104 57 109
rect 68 104 74 109
rect 85 104 91 109
rect 122 104 128 109
rect 143 104 149 109
rect 166 104 172 109
rect 177 104 183 109
rect 194 104 200 109
rect 205 104 211 109
rect 228 104 234 109
rect 249 104 255 109
rect 266 104 272 109
rect 301 104 307 109
rect 318 104 324 109
rect 335 104 341 109
rect 367 104 373 109
rect 384 104 390 109
rect 19 65 25 70
rect 14 63 25 65
rect 14 57 16 63
rect 22 57 25 63
rect 14 55 25 57
rect 19 36 25 55
rect 51 52 57 70
rect 68 68 74 70
rect 85 68 91 70
rect 68 66 80 68
rect 68 60 70 66
rect 76 60 80 66
rect 68 58 80 60
rect 85 66 99 68
rect 85 60 90 66
rect 96 60 99 66
rect 122 65 128 70
rect 143 68 149 70
rect 136 66 149 68
rect 85 58 99 60
rect 120 63 131 65
rect 51 50 63 52
rect 51 44 55 50
rect 61 44 63 50
rect 51 42 63 44
rect 68 43 74 58
rect 85 43 91 58
rect 120 57 123 63
rect 129 57 131 63
rect 136 60 138 66
rect 144 65 149 66
rect 144 60 146 65
rect 166 60 172 70
rect 177 68 183 70
rect 194 68 200 70
rect 177 61 200 68
rect 205 61 211 70
rect 228 68 234 70
rect 228 66 240 68
rect 228 65 232 66
rect 136 58 146 60
rect 120 55 131 57
rect 151 55 172 60
rect 54 36 60 42
rect 68 38 77 43
rect 71 36 77 38
rect 82 39 91 43
rect 82 36 88 39
rect 122 36 128 55
rect 151 51 157 55
rect 139 49 157 51
rect 139 43 142 49
rect 148 43 157 49
rect 139 41 157 43
rect 162 48 172 50
rect 185 48 191 61
rect 205 56 225 61
rect 230 60 232 65
rect 238 60 240 66
rect 230 58 240 60
rect 249 57 255 70
rect 266 65 272 70
rect 266 63 276 65
rect 266 57 268 63
rect 274 57 276 63
rect 220 53 225 56
rect 247 55 257 57
rect 220 51 237 53
rect 162 43 164 48
rect 170 43 172 48
rect 162 41 172 43
rect 143 36 149 41
rect 166 36 172 41
rect 177 46 191 48
rect 205 49 215 51
rect 177 40 180 46
rect 186 40 200 46
rect 177 38 200 40
rect 177 36 183 38
rect 194 36 200 38
rect 205 44 207 49
rect 213 44 215 49
rect 220 46 228 51
rect 205 42 215 44
rect 226 45 228 46
rect 234 45 237 51
rect 247 49 249 55
rect 255 49 257 55
rect 247 47 257 49
rect 266 55 276 57
rect 226 43 237 45
rect 205 36 211 42
rect 228 36 234 43
rect 249 36 255 47
rect 266 36 272 55
rect 301 49 307 70
rect 291 47 307 49
rect 291 41 294 47
rect 300 46 307 47
rect 318 65 324 70
rect 318 63 328 65
rect 318 57 320 63
rect 326 57 328 63
rect 318 55 328 57
rect 300 41 310 46
rect 318 43 324 55
rect 335 50 341 70
rect 367 59 373 70
rect 384 67 390 70
rect 291 39 310 41
rect 304 36 310 39
rect 315 38 324 43
rect 330 48 341 50
rect 362 57 373 59
rect 379 65 390 67
rect 379 60 381 65
rect 386 60 390 65
rect 379 58 390 60
rect 362 51 364 57
rect 370 51 373 57
rect 362 49 373 51
rect 330 43 332 48
rect 338 43 341 48
rect 330 41 341 43
rect 315 36 321 38
rect 332 36 338 41
rect 367 36 373 49
rect 384 36 390 58
rect 19 14 25 19
rect 54 14 60 19
rect 71 14 77 19
rect 82 14 88 19
rect 122 14 128 19
rect 143 14 149 19
rect 166 14 172 19
rect 177 14 183 19
rect 194 14 200 19
rect 205 14 211 19
rect 228 14 234 19
rect 249 14 255 19
rect 266 14 272 19
rect 304 14 310 19
rect 315 14 321 19
rect 332 14 338 19
rect 367 14 373 19
rect 384 14 390 19
<< polycontact >>
rect 16 57 22 63
rect 70 60 76 66
rect 90 60 96 66
rect 55 44 61 50
rect 123 57 129 63
rect 138 60 144 66
rect 142 43 148 49
rect 232 60 238 66
rect 268 57 274 63
rect 164 43 170 48
rect 180 40 186 46
rect 207 44 213 49
rect 228 45 234 51
rect 249 49 255 55
rect 294 41 300 47
rect 320 57 326 63
rect 381 60 386 65
rect 364 51 370 57
rect 332 43 338 48
<< metal1 >>
rect 0 118 410 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 131 118
rect 137 112 155 118
rect 161 112 179 118
rect 185 112 203 118
rect 209 112 227 118
rect 233 112 251 118
rect 257 112 275 118
rect 281 112 299 118
rect 305 112 323 118
rect 329 112 347 118
rect 353 112 371 118
rect 377 112 410 118
rect 0 111 410 112
rect 11 102 16 111
rect 11 70 16 72
rect 28 102 33 104
rect 16 63 22 65
rect 16 55 22 57
rect 28 51 33 72
rect 43 102 48 104
rect 28 50 34 51
rect 34 44 36 50
rect 28 38 34 44
rect 43 38 48 88
rect 60 102 65 104
rect 60 80 65 87
rect 77 102 82 111
rect 77 85 82 87
rect 94 102 99 104
rect 114 102 119 111
rect 114 95 119 97
rect 152 102 163 104
rect 94 80 99 87
rect 60 75 99 80
rect 108 86 152 90
rect 108 84 163 86
rect 186 102 191 111
rect 108 66 114 84
rect 186 82 191 84
rect 214 102 225 104
rect 258 102 263 111
rect 258 95 263 97
rect 275 102 280 104
rect 247 84 249 90
rect 255 84 257 90
rect 249 82 255 84
rect 220 74 225 76
rect 293 102 298 104
rect 293 80 298 87
rect 310 102 315 111
rect 310 85 315 87
rect 327 102 332 104
rect 327 80 332 87
rect 280 74 286 77
rect 293 75 332 80
rect 344 102 349 104
rect 344 82 349 88
rect 359 102 364 104
rect 344 77 350 82
rect 214 71 220 73
rect 275 72 286 74
rect 68 60 70 66
rect 76 60 78 66
rect 88 60 90 66
rect 96 60 114 66
rect 108 50 114 60
rect 121 57 123 63
rect 129 57 131 63
rect 136 60 138 66
rect 144 60 232 66
rect 238 63 274 66
rect 238 60 268 63
rect 53 44 55 50
rect 61 44 63 50
rect 108 44 131 50
rect 164 49 170 60
rect 207 49 213 60
rect 266 57 268 60
rect 274 57 276 63
rect 228 51 234 54
rect 77 38 95 44
rect 101 38 103 44
rect 11 34 16 36
rect 11 12 16 21
rect 28 34 33 38
rect 43 33 82 38
rect 63 32 82 33
rect 125 33 131 44
rect 140 43 142 49
rect 148 43 150 49
rect 162 48 172 49
rect 162 43 164 48
rect 170 43 172 48
rect 180 46 186 47
rect 178 40 180 46
rect 186 40 188 46
rect 205 44 207 49
rect 213 44 215 49
rect 247 49 249 55
rect 255 49 257 55
rect 281 50 286 72
rect 291 57 293 63
rect 299 57 313 63
rect 318 57 320 63
rect 326 57 328 63
rect 345 57 350 77
rect 376 102 381 111
rect 393 102 398 104
rect 376 81 381 83
rect 392 89 393 91
rect 392 81 393 83
rect 364 73 380 76
rect 359 70 380 73
rect 386 70 388 76
rect 380 69 386 70
rect 381 65 386 69
rect 228 44 234 45
rect 275 44 286 50
rect 228 39 280 44
rect 292 41 294 47
rect 300 41 302 47
rect 214 37 220 39
rect 63 31 68 32
rect 28 19 33 21
rect 46 26 51 28
rect 46 12 51 21
rect 63 19 68 21
rect 91 27 96 29
rect 91 12 96 21
rect 114 27 119 30
rect 125 28 163 33
rect 275 34 280 39
rect 307 38 313 57
rect 345 51 364 57
rect 370 51 372 57
rect 330 43 332 49
rect 338 43 340 49
rect 345 38 350 51
rect 381 42 386 60
rect 220 31 225 33
rect 114 12 119 21
rect 152 27 163 28
rect 152 19 163 21
rect 186 26 191 28
rect 186 12 191 21
rect 214 26 225 31
rect 214 19 225 21
rect 258 31 263 34
rect 258 12 263 21
rect 275 19 280 21
rect 296 34 301 36
rect 307 33 350 38
rect 359 37 386 42
rect 359 34 364 37
rect 296 12 301 21
rect 324 29 329 33
rect 324 19 329 21
rect 341 26 346 28
rect 341 12 346 21
rect 393 34 398 72
rect 359 19 364 21
rect 376 30 381 32
rect 376 12 381 21
rect 393 19 398 21
rect 0 11 410 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 131 11
rect 137 5 155 11
rect 161 5 179 11
rect 185 5 203 11
rect 209 5 227 11
rect 233 5 251 11
rect 257 5 275 11
rect 281 5 299 11
rect 305 5 323 11
rect 329 5 347 11
rect 353 5 371 11
rect 377 5 410 11
rect 0 0 410 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 36 118
rect 36 113 41 118
rect 35 112 41 113
rect 59 113 60 118
rect 60 113 65 118
rect 59 112 65 113
rect 83 113 84 118
rect 84 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 131 113 136 118
rect 136 113 137 118
rect 131 112 137 113
rect 155 113 160 118
rect 160 113 161 118
rect 155 112 161 113
rect 179 113 184 118
rect 184 113 185 118
rect 179 112 185 113
rect 203 113 208 118
rect 208 113 209 118
rect 203 112 209 113
rect 227 113 232 118
rect 232 113 233 118
rect 227 112 233 113
rect 251 113 256 118
rect 256 113 257 118
rect 251 112 257 113
rect 275 113 280 118
rect 280 113 281 118
rect 275 112 281 113
rect 299 113 304 118
rect 304 113 305 118
rect 299 112 305 113
rect 323 113 328 118
rect 328 113 329 118
rect 323 112 329 113
rect 347 113 352 118
rect 352 113 353 118
rect 347 112 353 113
rect 371 113 376 118
rect 376 113 377 118
rect 371 112 377 113
rect 16 57 22 63
rect 28 44 34 50
rect 249 84 255 90
rect 214 76 220 79
rect 214 73 220 76
rect 70 60 76 66
rect 90 60 96 66
rect 123 57 129 63
rect 55 44 61 50
rect 268 57 274 63
rect 95 38 101 44
rect 142 43 148 49
rect 180 40 186 46
rect 228 45 234 51
rect 249 49 255 55
rect 293 57 299 63
rect 320 57 326 63
rect 392 83 393 89
rect 393 83 398 89
rect 380 70 386 76
rect 294 41 300 47
rect 214 31 220 37
rect 364 51 370 57
rect 332 48 338 49
rect 332 43 338 48
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 36 10
rect 36 5 41 10
rect 59 10 65 11
rect 59 5 60 10
rect 60 5 65 10
rect 83 10 89 11
rect 83 5 84 10
rect 84 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 131 10 137 11
rect 131 5 136 10
rect 136 5 137 10
rect 155 10 161 11
rect 155 5 160 10
rect 160 5 161 10
rect 179 10 185 11
rect 179 5 184 10
rect 184 5 185 10
rect 203 10 209 11
rect 203 5 208 10
rect 208 5 209 10
rect 227 10 233 11
rect 227 5 232 10
rect 232 5 233 10
rect 251 10 257 11
rect 251 5 256 10
rect 256 5 257 10
rect 275 10 281 11
rect 275 5 280 10
rect 280 5 281 10
rect 299 10 305 11
rect 299 5 304 10
rect 304 5 305 10
rect 323 10 329 11
rect 323 5 328 10
rect 328 5 329 10
rect 347 10 353 11
rect 347 5 352 10
rect 352 5 353 10
rect 371 10 377 11
rect 371 5 376 10
rect 376 5 377 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 274 118 282 119
rect 298 118 306 119
rect 322 118 330 119
rect 346 118 354 119
rect 370 118 378 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 129 112 131 118
rect 137 112 139 118
rect 153 112 155 118
rect 161 112 163 118
rect 177 112 179 118
rect 185 112 187 118
rect 201 112 203 118
rect 209 112 211 118
rect 225 112 227 118
rect 233 112 235 118
rect 249 112 251 118
rect 257 112 259 118
rect 273 112 275 118
rect 281 112 283 118
rect 297 112 299 118
rect 305 112 307 118
rect 321 112 323 118
rect 329 112 331 118
rect 345 112 347 118
rect 353 112 355 118
rect 369 112 371 118
rect 377 112 379 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 274 111 282 112
rect 298 111 306 112
rect 322 111 330 112
rect 346 111 354 112
rect 370 111 378 112
rect 70 99 326 105
rect 70 67 76 99
rect 142 87 234 93
rect 248 90 256 91
rect 68 66 78 67
rect 15 63 23 64
rect 14 57 16 63
rect 22 57 24 63
rect 68 60 70 66
rect 76 60 78 66
rect 68 59 78 60
rect 88 66 98 67
rect 88 60 90 66
rect 96 60 98 66
rect 121 63 131 64
rect 88 59 98 60
rect 120 57 123 63
rect 129 57 132 63
rect 15 56 23 57
rect 121 56 131 57
rect 27 50 35 51
rect 53 50 63 51
rect 142 50 148 87
rect 214 80 220 81
rect 213 79 221 80
rect 213 73 214 79
rect 220 73 221 79
rect 213 72 221 73
rect 26 44 28 50
rect 34 44 55 50
rect 61 44 63 50
rect 141 49 150 50
rect 27 43 35 44
rect 53 43 63 44
rect 93 44 103 45
rect 55 24 61 43
rect 93 38 95 44
rect 101 38 132 44
rect 140 43 142 49
rect 148 43 150 49
rect 180 47 186 48
rect 141 42 150 43
rect 179 46 187 47
rect 93 37 103 38
rect 126 36 132 38
rect 179 40 180 46
rect 186 40 188 46
rect 179 39 187 40
rect 179 36 186 39
rect 214 38 220 72
rect 228 52 234 87
rect 247 84 249 90
rect 255 84 290 90
rect 248 83 256 84
rect 249 56 255 83
rect 284 64 290 84
rect 320 64 326 99
rect 391 89 399 90
rect 390 83 392 89
rect 398 83 400 89
rect 391 82 399 83
rect 379 76 387 77
rect 378 70 380 76
rect 386 70 388 76
rect 379 69 387 70
rect 267 63 275 64
rect 284 63 301 64
rect 266 57 268 63
rect 274 57 276 63
rect 284 57 293 63
rect 299 57 301 63
rect 267 56 275 57
rect 291 56 301 57
rect 318 63 328 64
rect 318 57 320 63
rect 326 57 328 63
rect 363 57 371 58
rect 318 56 328 57
rect 248 55 256 56
rect 227 51 235 52
rect 227 45 228 51
rect 234 45 235 51
rect 247 49 249 55
rect 255 49 257 55
rect 360 51 364 57
rect 370 51 372 57
rect 332 50 338 51
rect 363 50 371 51
rect 331 49 339 50
rect 248 48 256 49
rect 227 44 235 45
rect 292 47 302 48
rect 228 43 234 44
rect 292 41 294 47
rect 300 41 302 47
rect 292 40 302 41
rect 331 43 332 49
rect 338 43 339 49
rect 331 41 339 43
rect 213 37 221 38
rect 292 37 300 40
rect 126 30 186 36
rect 212 31 214 37
rect 220 31 300 37
rect 213 30 221 31
rect 331 24 337 41
rect 55 18 337 24
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 274 11 282 12
rect 298 11 306 12
rect 322 11 330 12
rect 346 11 354 12
rect 370 11 378 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 129 5 131 11
rect 137 5 139 11
rect 153 5 155 11
rect 161 5 163 11
rect 177 5 179 11
rect 185 5 187 11
rect 201 5 203 11
rect 209 5 211 11
rect 225 5 227 11
rect 233 5 235 11
rect 249 5 251 11
rect 257 5 259 11
rect 273 5 275 11
rect 281 5 283 11
rect 297 5 299 11
rect 305 5 307 11
rect 321 5 323 11
rect 329 5 331 11
rect 345 5 347 11
rect 353 5 355 11
rect 369 5 371 11
rect 377 5 379 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
rect 274 4 282 5
rect 298 4 306 5
rect 322 4 330 5
rect 346 4 354 5
rect 370 4 378 5
<< labels >>
rlabel metal2 13 8 13 8 1 GND
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 126 60 126 60 1 D
port 1 n
rlabel metal2 271 60 271 60 1 CLK
port 6 n
rlabel metal2 323 60 323 60 1 SN
port 8 n
rlabel metal2 395 86 395 86 1 Q
port 4 n
rlabel metal2 383 73 383 73 1 QN
port 5 n
rlabel metal2 19 60 19 60 1 RN
port 7 n
<< end >>
