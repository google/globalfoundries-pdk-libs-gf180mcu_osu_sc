magic
tech gf180mcuC
timestamp 1661532203
<< nwell >>
rect 0 97 62 159
<< nmos >>
rect 22 55 28 72
rect 33 55 39 72
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
<< ndiff >>
rect 12 63 22 72
rect 12 57 14 63
rect 19 57 22 63
rect 12 55 22 57
rect 28 55 33 72
rect 39 70 49 72
rect 39 57 42 70
rect 47 57 49 70
rect 39 55 49 57
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 113 28 138
rect 33 113 36 138
rect 25 106 36 113
rect 42 138 52 140
rect 42 108 45 138
rect 50 108 52 138
rect 42 106 52 108
<< ndiffc >>
rect 14 57 19 63
rect 42 57 47 70
<< pdiffc >>
rect 11 108 16 138
rect 28 113 33 138
rect 45 108 50 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 19 88 25 106
rect 11 86 25 88
rect 11 80 14 86
rect 20 80 25 86
rect 11 78 25 80
rect 19 77 25 78
rect 36 101 42 106
rect 36 99 50 101
rect 36 93 42 99
rect 48 93 50 99
rect 36 91 50 93
rect 36 77 42 91
rect 19 74 28 77
rect 22 72 28 74
rect 33 74 42 77
rect 33 72 39 74
rect 22 50 28 55
rect 33 50 39 55
<< polycontact >>
rect 14 80 20 86
rect 42 93 48 99
<< metal1 >>
rect 0 154 62 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 62 154
rect 0 147 62 148
rect 11 138 16 147
rect 28 138 33 140
rect 28 112 33 113
rect 45 138 50 147
rect 11 106 16 108
rect 26 106 28 112
rect 34 106 36 112
rect 45 106 50 108
rect 12 80 14 86
rect 20 80 22 86
rect 28 71 33 106
rect 40 93 42 99
rect 48 93 50 99
rect 14 66 33 71
rect 42 70 47 72
rect 14 63 19 66
rect 14 55 19 57
rect 42 48 47 57
rect 0 47 62 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 62 47
rect 0 36 62 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 28 106 34 112
rect 14 80 20 86
rect 42 93 48 99
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 10 147 18 148
rect 34 147 42 148
rect 26 112 36 113
rect 26 106 28 112
rect 34 106 36 112
rect 26 105 36 106
rect 40 99 50 100
rect 40 93 42 99
rect 48 93 50 99
rect 40 92 50 93
rect 12 86 22 87
rect 12 80 14 86
rect 20 80 22 86
rect 12 79 22 80
rect 10 47 18 48
rect 34 47 42 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 10 40 18 41
rect 34 40 42 41
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 14 44 14 44 1 GND
rlabel metal2 17 83 17 83 1 A
port 1 n
rlabel metal2 31 109 31 109 1 Y
port 3 n
rlabel metal2 45 96 45 96 1 B
port 2 n
<< end >>
