* NGSPICE file created from sky130_fd_pr__rf_pnp_05v5_W3p40L3p40.ext - technology: sky130A

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5 area=1.81611e+13p
.ends

