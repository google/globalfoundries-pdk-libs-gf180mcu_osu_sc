* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1__generic_slope = 0.0
* statistics {
*   mismatch {
*     vary  sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1__generic_slope dist=gauss std=1.0
*   }
* }
.include "sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_01p8x01p8_m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_shieldl1.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_shieldl1.model.spice"
.include "sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_shieldl1.model.spice"
.include "sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_shieldpo_floatm3.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_shieldpo_floatm3.model.spice"
.include "sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2_shieldpom3.model.spice"
.include "sky130_fd_pr__cap_vpp_03p9x03p9_m1m2_shieldl1_floatm3.model.spice"
.include "sky130_fd_pr__cap_vpp_08p6x07p8_l1m1m2_noshield_o1.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_l1m1m2_noshield_o1.model.spice"
.include "sky130_fd_pr__cap_vpp_08p6x07p8_m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2.model.spice"
.include "sky130_fd_pr__cap_vpp_02p4x04p6_m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield.model.spice"
.include "sky130_fd_pr__cap_vpp_11p5x11p7_m1m2_noshield.model.spice"
