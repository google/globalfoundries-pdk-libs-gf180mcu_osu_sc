# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffn_1 0 0 ;
  SIZE 14.25 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 14.25 8.3 ;
        RECT 12.55 5.55 12.8 8.3 ;
        RECT 9.95 5.55 10.35 8.3 ;
        RECT 7.25 6.3 7.5 8.3 ;
        RECT 4.45 5.55 4.7 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14.25 0.7 ;
        RECT 12.55 0 12.8 1.9 ;
        RECT 9.95 0 10.35 1.55 ;
        RECT 7.25 0 7.5 1.9 ;
        RECT 4.45 0 4.7 1.5 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 9.5 2.95 10 3.25 ;
        RECT 9.6 2.85 9.9 3.35 ;
      LAYER Metal2 ;
        RECT 9.5 2.95 10 3.25 ;
        RECT 9.55 2.9 9.95 3.3 ;
      LAYER Via1 ;
        RECT 9.62 2.97 9.88 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 3.6 2.4 3.9 ;
      LAYER Metal2 ;
        RECT 1.75 3.6 2.55 3.9 ;
        RECT 1.9 3.55 2.4 3.95 ;
      LAYER Via1 ;
        RECT 2.02 3.62 2.28 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.4 4.9 13.9 5.25 ;
        RECT 13.4 4.85 13.85 5.25 ;
        RECT 13.4 1.05 13.65 7.25 ;
      LAYER Metal2 ;
        RECT 13.4 4.9 13.9 5.2 ;
        RECT 13.45 4.85 13.85 5.25 ;
      LAYER Via1 ;
        RECT 13.52 4.92 13.78 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.7 4.25 13.15 4.55 ;
        RECT 12.8 2.15 13.05 4.55 ;
        RECT 11.7 2.15 13.05 2.4 ;
        RECT 11.7 4.25 11.95 7.25 ;
        RECT 11.7 1.05 11.95 2.4 ;
      LAYER Metal2 ;
        RECT 12.65 4.25 13.15 4.55 ;
        RECT 12.7 4.2 13.1 4.6 ;
      LAYER Via1 ;
        RECT 12.77 4.27 13.03 4.53 ;
    END
  END QN
  OBS
    LAYER Metal2 ;
      RECT 6.75 4.85 7.15 5.25 ;
      RECT 6.7 4.9 11.15 5.2 ;
      RECT 10.85 2.95 11.15 5.2 ;
      RECT 11.95 2.9 12.35 3.3 ;
      RECT 10.85 2.95 12.4 3.25 ;
      RECT 10.25 1.75 10.65 2.15 ;
      RECT 9.5 1.8 10.7 2.1 ;
      RECT 5.8 1.6 6.2 2 ;
      RECT 5.75 1.65 9.9 1.95 ;
      RECT 5.75 1.75 10.65 1.95 ;
      RECT 8.9 4.2 9.3 4.6 ;
      RECT 7.7 4.2 8.1 4.6 ;
      RECT 6.05 4.2 6.55 4.6 ;
      RECT 3.25 4.2 3.7 4.6 ;
      RECT 3.25 4.25 9.35 4.55 ;
      RECT 8.05 2.9 8.45 3.3 ;
      RECT 6.1 2.9 6.5 3.3 ;
      RECT 6.05 2.95 8.55 3.25 ;
      RECT 6.8 3.55 7.2 3.95 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 4.1 2.25 4.5 2.65 ;
      RECT 0.45 2.25 0.85 2.65 ;
      RECT 0.4 2.3 4.55 2.6 ;
    LAYER Via1 ;
      RECT 12.02 2.97 12.28 3.23 ;
      RECT 10.32 1.82 10.58 2.08 ;
      RECT 8.97 4.27 9.23 4.53 ;
      RECT 8.12 2.97 8.38 3.23 ;
      RECT 7.77 4.27 8.03 4.53 ;
      RECT 6.87 3.62 7.13 3.88 ;
      RECT 6.82 4.92 7.08 5.18 ;
      RECT 6.17 2.97 6.43 3.23 ;
      RECT 6.17 4.27 6.43 4.53 ;
      RECT 5.87 1.67 6.13 1.93 ;
      RECT 4.17 2.32 4.43 2.58 ;
      RECT 3.37 4.27 3.63 4.53 ;
      RECT 0.52 2.32 0.78 2.58 ;
    LAYER Metal1 ;
      RECT 10.95 1.05 11.2 7.25 ;
      RECT 10.95 2.95 12.4 3.25 ;
      RECT 10.3 1.8 10.6 5.3 ;
      RECT 10.2 4.9 10.7 5.2 ;
      RECT 10.2 1.8 10.7 2.1 ;
      RECT 9.1 5.55 9.35 7.25 ;
      RECT 8.95 1.7 9.25 5.8 ;
      RECT 9.1 1.05 9.35 1.95 ;
      RECT 8.1 4.85 8.35 7.25 ;
      RECT 8.1 4.85 8.7 5.1 ;
      RECT 8.4 3.65 8.7 5.1 ;
      RECT 8.1 2.85 8.4 3.9 ;
      RECT 8.1 1.05 8.35 3.9 ;
      RECT 6.7 4.9 7.2 5.2 ;
      RECT 6.8 3.6 7.1 5.2 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 5.5 4.25 6.55 4.55 ;
      RECT 5.5 2.25 5.8 4.55 ;
      RECT 5.4 2.25 5.9 2.55 ;
      RECT 5.85 6.05 6.1 7.25 ;
      RECT 4.95 6.05 6.1 6.3 ;
      RECT 4.95 3.55 5.2 6.3 ;
      RECT 4.9 1.7 5.15 3.8 ;
      RECT 4.9 1.7 6.25 1.95 ;
      RECT 5.85 1.65 6.25 1.95 ;
      RECT 5.85 1.05 6.1 1.95 ;
      RECT 4.05 4.9 4.55 5.2 ;
      RECT 4.15 2.3 4.45 5.2 ;
      RECT 4.05 2.3 4.55 2.6 ;
      RECT 2.6 4.25 3.75 4.55 ;
      RECT 3.35 2.3 3.65 4.55 ;
      RECT 3.25 2.3 3.75 2.6 ;
      RECT 3.05 5.05 3.3 7.25 ;
      RECT 1.4 5.05 3.3 5.3 ;
      RECT 1.4 2.35 1.65 5.3 ;
      RECT 1.05 4.25 1.65 4.55 ;
      RECT 1.4 2.35 2.4 2.6 ;
      RECT 2 1.65 2.4 2.6 ;
      RECT 2 1.65 3.3 1.9 ;
      RECT 3.05 1.05 3.3 1.9 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.5 2.2 0.8 2.7 ;
      RECT 7.65 4.25 8.15 4.55 ;
      RECT 6.05 2.95 6.55 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffn_1
