# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dlatn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlatn_1 0 0 ;
  SIZE 11.3 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 11.3 6.15 ;
        RECT 9.6 4.2 9.85 6.15 ;
        RECT 8 3.55 8.25 6.15 ;
        RECT 5.35 3.75 5.6 6.15 ;
        RECT 1.45 4.3 1.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 11.3 0.6 ;
        RECT 9.6 0 9.85 1.45 ;
        RECT 8 0 8.25 1.8 ;
        RECT 5.2 0 5.6 1.45 ;
        RECT 1.45 0 1.85 1.5 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.75 2.85 8.25 3.15 ;
      LAYER MET2 ;
        RECT 7.75 2.8 8.25 3.2 ;
      LAYER VIA12 ;
        RECT 7.87 2.87 8.13 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.45 2.85 10.95 3.15 ;
        RECT 10.45 2.8 10.85 3.2 ;
        RECT 10.45 0.95 10.7 5.2 ;
      LAYER MET2 ;
        RECT 10.45 2.85 10.95 3.15 ;
        RECT 10.5 2.8 10.9 3.2 ;
      LAYER VIA12 ;
        RECT 10.57 2.87 10.83 3.13 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 9 2.3 9.5 2.7 ;
      RECT 5.05 2.3 5.5 2.7 ;
      RECT 8.95 2.3 9.5 2.65 ;
      RECT 4.6 2.3 5.5 2.65 ;
      RECT 0.35 2.15 0.85 2.55 ;
      RECT 0.35 2.2 4.9 2.5 ;
      RECT 5.2 2.15 9.25 2.45 ;
      RECT 6.95 2.95 7.45 3.35 ;
      RECT 5.7 2.95 6.2 3.35 ;
      RECT 3.5 3 7.45 3.3 ;
      RECT 3.45 2.8 3.85 3.2 ;
      RECT 3.4 2.85 3.9 3.15 ;
    LAYER VIA12 ;
      RECT 9.12 2.37 9.38 2.63 ;
      RECT 7.07 3.02 7.33 3.28 ;
      RECT 5.82 3.02 6.08 3.28 ;
      RECT 5.12 2.37 5.38 2.63 ;
      RECT 3.52 2.87 3.78 3.13 ;
      RECT 0.47 2.22 0.73 2.48 ;
    LAYER MET1 ;
      RECT 8.75 3.35 9 5.2 ;
      RECT 8.75 3.35 10.1 3.6 ;
      RECT 9.8 1.85 10.1 3.6 ;
      RECT 8.75 1.85 10.1 2.1 ;
      RECT 8.75 0.95 9 2.1 ;
      RECT 7.15 0.95 7.4 5.2 ;
      RECT 6.95 3 7.45 3.3 ;
      RECT 6.2 3.65 6.45 5.2 ;
      RECT 6.45 2 6.7 3.9 ;
      RECT 2.6 3 3.1 3.3 ;
      RECT 2.7 2.3 3 3.3 ;
      RECT 4.15 2.45 4.65 2.75 ;
      RECT 2.7 2.3 4.5 2.6 ;
      RECT 2.7 2.35 4.55 2.6 ;
      RECT 4.2 1.7 4.5 2.75 ;
      RECT 6.2 0.95 6.45 2.25 ;
      RECT 4.2 1.7 6.45 1.95 ;
      RECT 3.15 3.8 3.4 5.2 ;
      RECT 1.15 3.8 3.4 4.05 ;
      RECT 1.15 1.9 1.4 4.05 ;
      RECT 1.1 3 1.55 3.3 ;
      RECT 1.15 1.9 2.4 2.15 ;
      RECT 2.15 1.2 2.4 2.15 ;
      RECT 3.15 0.95 3.4 1.55 ;
      RECT 2.15 1.2 3.4 1.45 ;
      RECT 0.6 0.95 0.85 5.2 ;
      RECT 0.5 2.15 0.85 2.55 ;
      RECT 0.35 2.2 0.85 2.5 ;
      RECT 0.45 2.15 0.85 2.5 ;
      RECT 9 2.35 9.5 2.65 ;
      RECT 5.7 3 6.2 3.3 ;
      RECT 5 2.35 5.5 2.65 ;
      RECT 3.4 2.85 3.9 3.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlatn_1
