* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__dlatn_1 D Q CLKN
X0 a_52_92 CLKN VDD VDD pmos_3p3 w=34 l=6
X1 a_46_19 D VSS VSS nmos_3p3 w=17 l=6
X2 a_20_14 CLKN a_46_19 VSS nmos_3p3 w=17 l=6
X3 VSS a_10_19 a_127_19 VSS nmos_3p3 w=17 l=6
X4 VDD a_10_19 a_77_109 VDD pmos_3p3 w=34 l=6
X5 a_77_109 CLKN a_20_14 VDD pmos_3p3 w=34 l=6
X6 a_20_14 a_52_92 a_43_109 VDD pmos_3p3 w=34 l=6
X7 VDD a_20_14 a_10_19 VDD pmos_3p3 w=34 l=6
X8 a_43_109 D VDD VDD pmos_3p3 w=34 l=6
X9 Q a_127_19 VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_10_19 a_127_19 VDD pmos_3p3 w=34 l=6
X11 a_77_19 a_52_92 a_20_14 VSS nmos_3p3 w=17 l=6
X12 Q a_127_19 VSS VSS nmos_3p3 w=17 l=6
X13 VSS a_10_19 a_77_19 VSS nmos_3p3 w=17 l=6
X14 a_52_92 CLKN VSS VSS nmos_3p3 w=17 l=6
X15 VSS a_20_14 a_10_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
