* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dffsr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dffsr_1 D Q QN SN RN CLK VDD VSS
X0 VSS a_41_72# a_172_21# VSS nfet_03p3 w=0.85u l=0.3u
X1 a_128_72# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 VDD a_247_49# QN VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS a_247_49# a_234_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VDD SN a_57_72# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_291_72# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_57_72# a_25_21# a_41_72# VDD pfet_03p3 w=1.7u l=0.3u
X8 a_200_72# a_41_72# VDD VDD pfet_03p3 w=1.7u l=0.3u
X9 VDD a_211_21# a_291_72# VDD pfet_03p3 w=1.7u l=0.3u
X10 a_41_72# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 a_128_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_247_49# QN VSS nfet_03p3 w=0.85u l=0.3u
X13 a_310_21# a_211_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 a_211_21# a_139_43# a_200_72# VDD pfet_03p3 w=1.7u l=0.3u
X15 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 a_139_43# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X17 a_82_16# CLK a_128_72# VDD pfet_03p3 w=1.7u l=0.3u
X18 a_200_21# a_41_72# VSS VSS nfet_03p3 w=0.85u l=0.3u
X19 a_247_49# SN a_310_21# VSS nfet_03p3 w=0.85u l=0.3u
X20 a_211_21# CLK a_200_21# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_57_72# a_82_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X23 a_82_16# a_139_43# a_128_21# VSS nfet_03p3 w=0.85u l=0.3u
X24 a_139_43# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 a_234_72# CLK a_211_21# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_247_49# a_25_21# a_291_72# VDD pfet_03p3 w=1.7u l=0.3u
X27 a_172_72# a_139_43# a_82_16# VDD pfet_03p3 w=1.7u l=0.3u
X28 a_77_21# SN a_41_72# VSS nfet_03p3 w=0.85u l=0.3u
X29 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X30 VDD a_41_72# a_172_72# VDD pfet_03p3 w=1.7u l=0.3u
X31 a_234_21# a_139_43# a_211_21# VSS nfet_03p3 w=0.85u l=0.3u
X32 a_172_21# CLK a_82_16# VSS nfet_03p3 w=0.85u l=0.3u
X33 VSS a_82_16# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X34 VSS a_25_21# a_247_49# VSS nfet_03p3 w=0.85u l=0.3u
X35 VDD a_247_49# a_234_72# VDD pfet_03p3 w=1.7u l=0.3u
.ends
