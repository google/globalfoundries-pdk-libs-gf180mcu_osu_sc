* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_mux2_1 Y Sel A B
X0 B Sel Y VSS nmos_3p3 w=17 l=6
X1 Y a_23_16 A VSS nmos_3p3 w=17 l=6
X2 a_23_16 Sel VSS VSS nmos_3p3 w=17 l=6
X3 Y Sel A VDD pmos_3p3 w=34 l=6
X4 B a_23_16 Y VDD pmos_3p3 w=34 l=6
X5 a_23_16 Sel VDD VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
