# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_mux2_1
  CLASS CORE ;
  ORIGIN 0.1 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_mux2_1 -0.1 -0.15 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 3.3 2.75 3.7 ;
        RECT 2.15 0.8 2.4 7 ;
      LAYER MET2 ;
        RECT 2.25 3.3 2.75 3.7 ;
      LAYER VIA12 ;
        RECT 2.37 3.37 2.63 3.63 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.65 3.95 4.15 4.35 ;
        RECT 3.85 0.8 4.1 7 ;
      LAYER MET2 ;
        RECT 3.65 3.95 4.15 4.35 ;
      LAYER VIA12 ;
        RECT 3.77 4.02 4.03 4.28 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.7 0.95 3 ;
      LAYER MET2 ;
        RECT 0.45 2.65 0.95 3.05 ;
      LAYER VIA12 ;
        RECT 0.57 2.72 0.83 2.98 ;
    END
  END Sel
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -0.1 7.35 4.7 7.95 ;
        RECT 0.45 5.3 0.7 7.95 ;
      LAYER MET2 ;
        RECT 2.75 7.4 3.25 7.7 ;
        RECT 2.8 7.35 3.2 7.75 ;
        RECT 1.55 7.4 2.05 7.7 ;
        RECT 1.6 7.35 2 7.75 ;
        RECT 0.35 7.4 0.85 7.7 ;
        RECT 0.4 7.35 0.8 7.75 ;
      LAYER VIA12 ;
        RECT 0.47 7.42 0.73 7.68 ;
        RECT 1.67 7.42 1.93 7.68 ;
        RECT 2.87 7.42 3.13 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -0.1 -0.15 4.7 0.45 ;
        RECT 0.45 -0.15 0.7 1.65 ;
      LAYER MET2 ;
        RECT 2.75 0.1 3.25 0.4 ;
        RECT 2.8 0.05 3.2 0.45 ;
        RECT 1.55 0.1 2.05 0.4 ;
        RECT 1.6 0.05 2 0.45 ;
        RECT 0.35 0.1 0.85 0.4 ;
        RECT 0.4 0.05 0.8 0.45 ;
      LAYER VIA12 ;
        RECT 0.47 0.12 0.73 0.38 ;
        RECT 1.67 0.12 1.93 0.38 ;
        RECT 2.87 0.12 3.13 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 4.6 3.4 5 ;
        RECT 3 0.8 3.25 7 ;
      LAYER MET2 ;
        RECT 2.9 4.6 3.4 5 ;
      LAYER VIA12 ;
        RECT 3.02 4.67 3.28 4.93 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.3 0.8 1.55 7 ;
      RECT 1.3 4 1.9 4.3 ;
      RECT 1.3 2.05 1.9 2.35 ;
  END
END gf180mcu_osu_sc_12T_mux2_1
