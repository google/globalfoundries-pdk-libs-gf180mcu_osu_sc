magic
tech gf180mcuC
timestamp 1661527449
<< nwell >>
rect 0 97 82 159
<< nmos >>
rect 22 55 28 72
rect 33 55 39 72
rect 57 55 63 72
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 57 106 63 140
<< ndiff >>
rect 12 62 22 72
rect 12 57 14 62
rect 19 57 22 62
rect 12 55 22 57
rect 28 55 33 72
rect 39 70 57 72
rect 39 57 42 70
rect 54 57 57 70
rect 39 55 57 57
rect 63 62 73 72
rect 63 57 66 62
rect 71 57 73 62
rect 63 55 73 57
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 108 28 138
rect 33 108 36 138
rect 25 106 36 108
rect 42 138 57 140
rect 42 108 45 138
rect 54 108 57 138
rect 42 106 57 108
rect 63 138 73 140
rect 63 128 66 138
rect 71 128 73 138
rect 63 106 73 128
<< ndiffc >>
rect 14 57 19 62
rect 42 57 54 70
rect 66 57 71 62
<< pdiffc >>
rect 11 108 16 138
rect 28 108 33 138
rect 45 108 54 138
rect 66 128 71 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
rect 57 46 66 48
rect 57 41 59 46
rect 64 41 66 46
rect 57 39 66 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
rect 59 41 64 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 57 140 63 145
rect 19 88 25 106
rect 36 101 42 106
rect 36 99 49 101
rect 36 97 41 99
rect 11 86 25 88
rect 11 80 14 86
rect 20 82 25 86
rect 33 93 41 97
rect 47 93 49 99
rect 33 91 49 93
rect 20 80 28 82
rect 11 78 28 80
rect 22 72 28 78
rect 33 72 39 91
rect 57 88 63 106
rect 53 86 63 88
rect 53 80 55 86
rect 61 80 63 86
rect 53 78 63 80
rect 57 72 63 78
rect 22 50 28 55
rect 33 50 39 55
rect 57 50 63 55
<< polycontact >>
rect 14 80 20 86
rect 41 93 47 99
rect 55 80 61 86
<< metal1 >>
rect 0 154 82 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 82 154
rect 0 147 82 148
rect 11 138 16 147
rect 11 106 16 108
rect 28 138 33 140
rect 28 86 33 108
rect 45 138 54 147
rect 45 106 54 108
rect 66 138 71 140
rect 66 113 71 128
rect 66 112 74 113
rect 66 106 68 112
rect 74 106 76 112
rect 66 105 74 106
rect 39 93 41 99
rect 47 93 49 99
rect 55 86 61 88
rect 12 80 14 86
rect 20 80 22 86
rect 28 80 55 86
rect 28 70 33 80
rect 55 78 61 80
rect 14 65 33 70
rect 42 70 54 72
rect 14 62 19 65
rect 14 55 19 57
rect 42 48 54 57
rect 66 62 71 105
rect 66 55 71 57
rect 0 47 82 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 59 47
rect 65 41 82 47
rect 0 36 82 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 68 106 74 112
rect 41 93 47 99
rect 14 80 20 86
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
rect 59 46 65 47
rect 59 41 64 46
rect 64 41 65 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 66 112 76 113
rect 66 106 68 112
rect 74 106 76 112
rect 66 105 76 106
rect 39 99 49 100
rect 39 93 41 99
rect 47 93 49 99
rect 39 92 49 93
rect 13 86 21 87
rect 12 80 14 86
rect 20 80 22 86
rect 13 79 21 80
rect 10 47 18 48
rect 34 47 42 48
rect 58 47 66 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 57 41 59 47
rect 65 41 67 47
rect 10 40 18 41
rect 34 40 42 41
rect 58 40 66 41
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 17 83 17 83 1 A
port 1 n
rlabel metal2 14 44 14 44 1 GND
rlabel metal2 44 96 44 96 1 B
port 2 n
rlabel metal2 71 109 71 109 1 Y
port 3 n
<< end >>
