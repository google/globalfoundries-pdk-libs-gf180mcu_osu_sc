# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addh_1 0 0 ;
  SIZE 8.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 8.1 8.3 ;
        RECT 6.4 5.55 6.65 8.3 ;
        RECT 3.85 5.55 4.1 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 8.1 0.7 ;
        RECT 6.4 0 6.65 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.9 3.6 4.4 3.9 ;
        RECT 1.5 3.6 2 3.9 ;
      LAYER Metal2 ;
        RECT 3.9 3.55 4.4 3.95 ;
        RECT 1.5 3.6 4.4 3.9 ;
        RECT 1.5 3.55 2 3.95 ;
      LAYER Via1 ;
        RECT 1.62 3.62 1.88 3.88 ;
        RECT 4.02 3.62 4.28 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.2 2.95 5.7 3.25 ;
        RECT 2.35 2.95 2.85 3.25 ;
      LAYER Metal2 ;
        RECT 5.2 2.9 5.7 3.3 ;
        RECT 2.35 2.95 5.7 3.25 ;
        RECT 2.35 2.9 2.85 3.3 ;
      LAYER Via1 ;
        RECT 2.47 2.97 2.73 3.23 ;
        RECT 5.32 2.97 5.58 3.23 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 2.3 0.9 2.6 ;
        RECT 0.55 1.05 0.8 7.25 ;
      LAYER Metal2 ;
        RECT 0.4 2.25 0.9 2.65 ;
      LAYER Via1 ;
        RECT 0.52 2.32 0.78 2.58 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.2 4.9 7.7 5.2 ;
        RECT 7.25 4.85 7.6 5.25 ;
        RECT 7.25 1.05 7.5 7.25 ;
      LAYER Metal2 ;
        RECT 7.2 4.85 7.7 5.25 ;
      LAYER Via1 ;
        RECT 7.32 4.92 7.58 5.18 ;
    END
  END S
  OBS
    LAYER Metal2 ;
      RECT 6.05 4.85 6.55 5.25 ;
      RECT 3 4.85 3.5 5.25 ;
      RECT 3 4.9 6.55 5.2 ;
    LAYER Via1 ;
      RECT 6.17 4.92 6.43 5.18 ;
      RECT 3.12 4.92 3.38 5.18 ;
    LAYER Metal1 ;
      RECT 5.55 3.6 5.8 7.25 ;
      RECT 5.55 3.6 7 3.9 ;
      RECT 4.7 3.6 7 3.85 ;
      RECT 4.7 1.45 4.95 3.85 ;
      RECT 5.55 0.95 5.8 2 ;
      RECT 3.85 0.95 4.1 2 ;
      RECT 3.85 0.95 5.8 1.2 ;
      RECT 2.25 4.9 2.5 7.25 ;
      RECT 1.05 4.9 3.5 5.2 ;
      RECT 3.1 1.05 3.35 5.2 ;
      RECT 6.05 4.9 6.55 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addh_1
