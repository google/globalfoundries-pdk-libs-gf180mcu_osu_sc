* NGSPICE file created from gf180mcu_osu_sc_12T_addh_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 VDD B a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_19_14# CO VDD pmos_3p3 w=1.7u l=0.3u
X3 a_19_14# B a_42_19# GND nmos_3p3 w=0.85u l=0.3u
X4 S a_91_19# GND GND nmos_3p3 w=0.85u l=0.3u
X5 GND a_19_14# CO GND nmos_3p3 w=0.85u l=0.3u
X6 S a_91_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 a_91_19# B a_91_109# VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_19_14# a_91_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_91_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 a_91_19# A a_75_19# GND nmos_3p3 w=0.85u l=0.3u
X11 a_42_19# A GND GND nmos_3p3 w=0.85u l=0.3u
X12 GND a_19_14# a_75_19# GND nmos_3p3 w=0.85u l=0.3u
X13 a_75_19# B a_91_19# GND nmos_3p3 w=0.85u l=0.3u
