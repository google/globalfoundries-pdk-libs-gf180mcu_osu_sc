

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_tielo Y
X0 Y a_19_14 GND GND nmos_3p3 w=17 l=6
X1 a_19_14 a_19_14 VDD VDD pmos_3p3 w=34 l=6
.ends

