* SKY130 Spice File.
.include "../../sky130_fd_pr__nfet_01v8__fs.corner.spice"
.include "../../sky130_fd_pr__nfet_01v8__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_01v8_lvt__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_03v3_nvt__fs.corner.spice"
.include "../../sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_05v0_nvt__fs.corner.spice"
.include "../../sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__esd_nfet_01v8__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_lvt__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_lvt__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_hvt__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_hvt__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__esd_pfet_g5v0d10v5__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d10v5__fs.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d10v5__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d16v0__fs.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d10v5__fs.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d16v0__fs_discrete.corner.spice"
.include "../../sky130_fd_pr__esd_nfet_g5v0d10v5__fs.corner.spice"
.include "nonfet.spice"
.include "../../sky130_fd_pr__nfet_01v8_lvt__subvt_mismatch.corner.spice"
.include "../../sky130_fd_pr__pfet_20v0__fs_discrete.corner.spice"
.include "../../sky130_fd_pr__nfet_20v0__fs_discrete.corner.spice"
.include "../../sky130_fd_pr__nfet_20v0_nvt__fs_discrete.corner.spice"
.include "../../all.spice"
.include "rf.spice"
