* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__clkinv_16.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__clkinv_16 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X3 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X5 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X6 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X9 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X10 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X13 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X15 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X16 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X17 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X18 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X19 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X20 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X21 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X22 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X23 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X24 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X26 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X27 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X28 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X29 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X30 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
C0 Y VDD 2.062410fF
.ends
