# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dlat_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlat_1 0 0 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET2 ;
        RECT 5.2 4.1 5.7 4.5 ;
        RECT 3.45 4.15 5.7 4.45 ;
        RECT 3.5 4.1 3.9 4.5 ;
      LAYER MET1 ;
        RECT 5.2 4.15 5.7 4.45 ;
        RECT 3.45 4.15 3.95 4.45 ;
      LAYER VIA12 ;
        RECT 3.57 4.17 3.83 4.43 ;
        RECT 5.32 4.17 5.58 4.43 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 9 8.1 ;
        RECT 7.3 5.45 7.55 8.1 ;
        RECT 4.85 5.45 5.1 8.1 ;
        RECT 1.45 6.25 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9 0.6 ;
        RECT 7.3 0 7.55 1.8 ;
        RECT 4.7 0 5.1 1.8 ;
        RECT 1.45 0 1.85 1.8 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 1.85 4.1 2.35 4.5 ;
      LAYER MET1 ;
        RECT 1.85 4.15 2.35 4.45 ;
      LAYER VIA12 ;
        RECT 1.97 4.17 2.23 4.43 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 8.15 4.8 8.65 5.1 ;
        RECT 8.2 4.75 8.6 5.15 ;
      LAYER MET1 ;
        RECT 8.15 4.8 8.65 5.1 ;
        RECT 8.15 4.75 8.55 5.15 ;
        RECT 8.15 0.95 8.4 7.15 ;
      LAYER VIA12 ;
        RECT 8.27 4.82 8.53 5.08 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 6.75 3.45 7.25 3.85 ;
      RECT 4.55 3.45 4.95 3.85 ;
      RECT 0.35 3.45 0.85 3.85 ;
      RECT 0.35 3.5 7.25 3.8 ;
      RECT 6.5 4.75 6.9 5.15 ;
      RECT 6.45 4.8 6.95 5.1 ;
    LAYER VIA12 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.57 4.82 6.83 5.08 ;
      RECT 4.62 3.52 4.88 3.78 ;
      RECT 0.47 3.52 0.73 3.78 ;
    LAYER MET1 ;
      RECT 6.45 4.75 6.7 7.15 ;
      RECT 6.45 4.75 6.85 5.3 ;
      RECT 6.45 4.8 6.95 5.1 ;
      RECT 6.45 4.8 7.8 5.05 ;
      RECT 7.5 2.05 7.8 5.05 ;
      RECT 6.45 2.05 7.8 2.3 ;
      RECT 6.45 0.95 6.7 2.3 ;
      RECT 5.7 5.25 5.95 7.15 ;
      RECT 5.95 1.95 6.2 5.5 ;
      RECT 2.6 4.7 3.1 5 ;
      RECT 2.7 2.55 3 5 ;
      RECT 2.7 2.55 6.2 2.85 ;
      RECT 5.7 0.95 5.95 2.2 ;
      RECT 3.15 5.45 3.4 7.15 ;
      RECT 1.15 5.45 3.4 5.7 ;
      RECT 1.15 2.05 1.4 5.7 ;
      RECT 1.1 4.15 1.55 4.45 ;
      RECT 1.15 2.05 3.4 2.3 ;
      RECT 3.15 0.95 3.4 2.3 ;
      RECT 0.6 0.95 0.85 7.15 ;
      RECT 0.5 3.45 0.85 3.85 ;
      RECT 0.35 3.5 0.85 3.8 ;
      RECT 0.45 3.45 0.85 3.8 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.5 3.5 5 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlat_1
