# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dlatn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlatn_1 0 0 ;
  SIZE 11.3 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 11.3 6.35 ;
        RECT 9.6 4.3 9.85 6.35 ;
        RECT 8 3.65 8.25 6.35 ;
        RECT 5.35 3.85 5.6 6.35 ;
        RECT 1.45 4.4 1.7 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 11.3 0.7 ;
        RECT 9.6 0 9.85 1.55 ;
        RECT 8 0 8.25 1.9 ;
        RECT 5.2 0 5.6 1.55 ;
        RECT 1.45 0 1.85 1.6 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 7.75 2.95 8.25 3.25 ;
      LAYER Metal2 ;
        RECT 7.75 2.9 8.25 3.3 ;
      LAYER Via1 ;
        RECT 7.87 2.97 8.13 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.85 2.95 2.35 3.25 ;
      LAYER Metal2 ;
        RECT 1.85 2.9 2.35 3.3 ;
      LAYER Via1 ;
        RECT 1.97 2.97 2.23 3.23 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.45 2.95 10.95 3.25 ;
        RECT 10.45 2.9 10.85 3.3 ;
        RECT 10.45 1.05 10.7 5.3 ;
      LAYER Metal2 ;
        RECT 10.45 2.95 10.95 3.25 ;
        RECT 10.5 2.9 10.9 3.3 ;
      LAYER Via1 ;
        RECT 10.57 2.97 10.83 3.23 ;
    END
  END Q
  OBS
    LAYER Metal2 ;
      RECT 9 2.4 9.5 2.8 ;
      RECT 5.05 2.4 5.5 2.8 ;
      RECT 8.95 2.4 9.5 2.75 ;
      RECT 4.6 2.4 5.5 2.75 ;
      RECT 0.35 2.25 0.85 2.65 ;
      RECT 0.35 2.3 4.9 2.6 ;
      RECT 5.2 2.25 9.25 2.55 ;
      RECT 6.95 3.05 7.45 3.45 ;
      RECT 5.7 3.05 6.2 3.45 ;
      RECT 3.5 3.1 7.45 3.4 ;
      RECT 3.45 2.9 3.85 3.3 ;
      RECT 3.4 2.95 3.9 3.25 ;
    LAYER Via1 ;
      RECT 9.12 2.47 9.38 2.73 ;
      RECT 7.07 3.12 7.33 3.38 ;
      RECT 5.82 3.12 6.08 3.38 ;
      RECT 5.12 2.47 5.38 2.73 ;
      RECT 3.52 2.97 3.78 3.23 ;
      RECT 0.47 2.32 0.73 2.58 ;
    LAYER Metal1 ;
      RECT 8.75 3.45 9 5.3 ;
      RECT 8.75 3.45 10.1 3.7 ;
      RECT 9.8 1.95 10.1 3.7 ;
      RECT 8.75 1.95 10.1 2.2 ;
      RECT 8.75 1.05 9 2.2 ;
      RECT 7.15 1.05 7.4 5.3 ;
      RECT 6.95 3.1 7.45 3.4 ;
      RECT 6.2 3.75 6.45 5.3 ;
      RECT 6.45 2.1 6.7 4 ;
      RECT 2.6 3.1 3.1 3.4 ;
      RECT 2.7 2.4 3 3.4 ;
      RECT 4.15 2.55 4.65 2.85 ;
      RECT 2.7 2.4 4.5 2.7 ;
      RECT 2.7 2.45 4.55 2.7 ;
      RECT 4.2 1.8 4.5 2.85 ;
      RECT 6.2 1.05 6.45 2.35 ;
      RECT 4.2 1.8 6.45 2.05 ;
      RECT 3.15 3.9 3.4 5.3 ;
      RECT 1.15 3.9 3.4 4.15 ;
      RECT 1.15 2 1.4 4.15 ;
      RECT 1.1 3.1 1.55 3.4 ;
      RECT 1.15 2 2.4 2.25 ;
      RECT 2.15 1.3 2.4 2.25 ;
      RECT 3.15 1.05 3.4 1.65 ;
      RECT 2.15 1.3 3.4 1.55 ;
      RECT 0.6 1.05 0.85 5.3 ;
      RECT 0.5 2.25 0.85 2.65 ;
      RECT 0.35 2.3 0.85 2.6 ;
      RECT 0.45 2.25 0.85 2.6 ;
      RECT 9 2.45 9.5 2.75 ;
      RECT 5.7 3.1 6.2 3.4 ;
      RECT 5 2.45 5.5 2.75 ;
      RECT 3.4 2.95 3.9 3.4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlatn_1
