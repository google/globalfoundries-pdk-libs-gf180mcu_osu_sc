# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_clkinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_clkinv_4 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 4.45 3.35 4.7 ;
        RECT 2.95 4.35 3.35 4.7 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 2.95 4.35 3.45 4.75 ;
      LAYER VIA12 ;
        RECT 3.07 4.42 3.33 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_12T_clkinv_4
