# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__tbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tbuf_8 0 0 ;
  SIZE 9.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 9.8 8.1 ;
        RECT 8.95 5.45 9.2 8.1 ;
        RECT 7.25 5.45 7.5 8.1 ;
        RECT 5.55 5.45 5.8 8.1 ;
        RECT 3.85 5.45 4.1 8.1 ;
        RECT 2.15 5.45 2.4 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.8 0.6 ;
        RECT 8.95 0 9.2 1.8 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 2.15 0 2.4 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 4.15 2.3 4.45 ;
      LAYER MET2 ;
        RECT 1.8 4.15 2.3 4.45 ;
        RECT 1.85 4.1 2.25 4.5 ;
      LAYER VIA12 ;
        RECT 1.92 4.17 2.18 4.43 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 2.2 1.45 2.5 ;
      LAYER MET2 ;
        RECT 0.95 2.15 1.45 2.55 ;
      LAYER VIA12 ;
        RECT 1.07 2.22 1.33 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 4.8 1.45 5.1 ;
      LAYER MET2 ;
        RECT 0.95 4.75 1.45 5.15 ;
      LAYER VIA12 ;
        RECT 1.07 4.82 1.33 5.08 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8 4.8 8.5 5.1 ;
        RECT 8.1 0.95 8.35 7.15 ;
        RECT 3 4.85 8.35 5.15 ;
        RECT 3 2.05 8.35 2.3 ;
        RECT 6.4 0.95 6.65 7.15 ;
        RECT 4.7 0.95 4.95 7.15 ;
        RECT 3 0.95 3.25 7.15 ;
      LAYER MET2 ;
        RECT 7.95 4.85 8.5 5.15 ;
        RECT 8 4.75 8.5 5.15 ;
      LAYER VIA12 ;
        RECT 8.12 4.82 8.38 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.75 5.45 1 7.15 ;
      RECT 0.45 5.45 1 5.7 ;
      RECT 0.45 1.55 0.7 5.7 ;
      RECT 0.45 2.9 2.75 3.2 ;
      RECT 0.45 1.55 1 1.8 ;
      RECT 0.75 0.95 1 1.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tbuf_8
