* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_oai31_1 Y A0 A1 B A2
X0 a_25_19 A1 VSS VSS nmos_3p3 w=17 l=6
X1 a_25_19 A2 VSS VSS nmos_3p3 w=17 l=6
X2 Y A1 a_45_70 VDD pmos_3p3 w=34 l=6
X3 Y B a_25_19 VSS nmos_3p3 w=17 l=6
X4 a_34_70 A2 VDD VDD pmos_3p3 w=34 l=6
X5 VSS A0 a_25_19 VSS nmos_3p3 w=17 l=6
X6 a_45_70 A0 a_34_70 VDD pmos_3p3 w=34 l=6
X7 VDD B Y VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
