magic
tech gf180mcuC
timestamp 1661875083
<< nwell >>
rect 0 61 32 123
<< metal1 >>
rect 0 111 32 123
rect 0 0 32 12
<< labels >>
rlabel metal1 10 117 10 117 1 VDD
rlabel metal1 6 6 6 6 1 GND
<< end >>
