* NGSPICE file created from gf180mcu_osu_sc_9T_xor2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_42_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 GND a_52_59# a_81_19# GND nmos_3p3 w=0.85u l=0.3u
X2 VDD B a_81_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 Y B a_42_19# GND nmos_3p3 w=0.85u l=0.3u
X4 GND A a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X5 Y a_52_59# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_81_19# a_9_19# Y GND nmos_3p3 w=0.85u l=0.3u
X8 a_52_59# B GND GND nmos_3p3 w=0.85u l=0.3u
X9 a_81_70# a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X10 a_52_59# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X11 a_42_19# A GND GND nmos_3p3 w=0.85u l=0.3u
