magic
tech gf180mcuC
timestamp 1659647090
<< nwell >>
rect 0 100 280 162
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 53 19 59 36
rect 70 19 76 36
rect 87 19 93 36
rect 104 19 110 36
rect 121 19 127 36
rect 138 19 144 36
rect 155 19 161 36
rect 172 19 178 36
rect 189 19 195 36
rect 206 19 212 36
rect 223 19 229 36
rect 255 19 261 36
<< pmos >>
rect 19 109 25 143
rect 36 109 42 143
rect 53 109 59 143
rect 70 109 76 143
rect 87 109 93 143
rect 104 109 110 143
rect 121 109 127 143
rect 138 109 144 143
rect 155 109 161 143
rect 172 109 178 143
rect 189 109 195 143
rect 206 109 212 143
rect 223 109 229 143
rect 255 109 261 143
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 34 53 36
rect 42 21 45 34
rect 50 21 53 34
rect 42 19 53 21
rect 59 34 70 36
rect 59 21 62 34
rect 67 21 70 34
rect 59 19 70 21
rect 76 19 87 36
rect 93 34 104 36
rect 93 21 96 34
rect 101 21 104 34
rect 93 19 104 21
rect 110 33 121 36
rect 110 21 113 33
rect 118 21 121 33
rect 110 19 121 21
rect 127 27 138 36
rect 127 21 130 27
rect 135 21 138 27
rect 127 19 138 21
rect 144 33 155 36
rect 144 21 147 33
rect 152 21 155 33
rect 144 19 155 21
rect 161 34 172 36
rect 161 21 164 34
rect 169 21 172 34
rect 161 19 172 21
rect 178 19 189 36
rect 195 19 206 36
rect 212 34 223 36
rect 212 21 215 34
rect 220 21 223 34
rect 212 19 223 21
rect 229 34 239 36
rect 229 21 232 34
rect 237 21 239 34
rect 229 19 239 21
rect 245 34 255 36
rect 245 21 247 34
rect 252 21 255 34
rect 245 19 255 21
rect 261 34 271 36
rect 261 21 264 34
rect 269 21 271 34
rect 261 19 271 21
<< pdiff >>
rect 9 141 19 143
rect 9 111 11 141
rect 16 111 19 141
rect 9 109 19 111
rect 25 141 36 143
rect 25 111 28 141
rect 33 111 36 141
rect 25 109 36 111
rect 42 141 53 143
rect 42 111 45 141
rect 50 111 53 141
rect 42 109 53 111
rect 59 141 70 143
rect 59 111 62 141
rect 67 111 70 141
rect 59 109 70 111
rect 76 109 87 143
rect 93 141 104 143
rect 93 111 96 141
rect 101 111 104 141
rect 93 109 104 111
rect 110 141 121 143
rect 110 111 113 141
rect 118 111 121 141
rect 110 109 121 111
rect 127 141 138 143
rect 127 111 130 141
rect 135 111 138 141
rect 127 109 138 111
rect 144 141 155 143
rect 144 111 147 141
rect 152 111 155 141
rect 144 109 155 111
rect 161 141 172 143
rect 161 111 164 141
rect 169 111 172 141
rect 161 109 172 111
rect 178 109 189 143
rect 195 109 206 143
rect 212 141 223 143
rect 212 111 215 141
rect 220 111 223 141
rect 212 109 223 111
rect 229 141 239 143
rect 229 111 232 141
rect 237 111 239 141
rect 229 109 239 111
rect 245 141 255 143
rect 245 111 247 141
rect 252 111 255 141
rect 245 109 255 111
rect 261 141 271 143
rect 261 111 264 141
rect 269 111 271 141
rect 261 109 271 111
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 45 21 50 34
rect 62 21 67 34
rect 96 21 101 34
rect 113 21 118 33
rect 130 21 135 27
rect 147 21 152 33
rect 164 21 169 34
rect 215 21 220 34
rect 232 21 237 34
rect 247 21 252 34
rect 264 21 269 34
<< pdiffc >>
rect 11 111 16 141
rect 28 111 33 141
rect 45 111 50 141
rect 62 111 67 141
rect 96 111 101 141
rect 113 111 118 141
rect 130 111 135 141
rect 147 111 152 141
rect 164 111 169 141
rect 215 111 220 141
rect 232 111 237 141
rect 247 111 252 141
rect 264 111 269 141
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 129 10 138 12
rect 129 5 131 10
rect 136 5 138 10
rect 129 3 138 5
rect 153 10 162 12
rect 153 5 155 10
rect 160 5 162 10
rect 153 3 162 5
rect 177 10 186 12
rect 177 5 179 10
rect 184 5 186 10
rect 177 3 186 5
rect 201 10 210 12
rect 201 5 203 10
rect 208 5 210 10
rect 201 3 210 5
rect 225 10 234 12
rect 225 5 227 10
rect 232 5 234 10
rect 225 3 234 5
rect 249 10 258 12
rect 249 5 251 10
rect 256 5 258 10
rect 249 3 258 5
<< nsubdiff >>
rect 9 157 18 159
rect 9 152 11 157
rect 16 152 18 157
rect 9 150 18 152
rect 33 157 42 159
rect 33 152 35 157
rect 40 152 42 157
rect 33 150 42 152
rect 57 157 66 159
rect 57 152 59 157
rect 64 152 66 157
rect 57 150 66 152
rect 81 157 90 159
rect 81 152 83 157
rect 88 152 90 157
rect 81 150 90 152
rect 105 157 114 159
rect 105 152 107 157
rect 112 152 114 157
rect 105 150 114 152
rect 129 157 138 159
rect 129 152 131 157
rect 136 152 138 157
rect 129 150 138 152
rect 153 157 162 159
rect 153 152 155 157
rect 160 152 162 157
rect 153 150 162 152
rect 177 157 186 159
rect 177 152 179 157
rect 184 152 186 157
rect 177 150 186 152
rect 201 157 210 159
rect 201 152 203 157
rect 208 152 210 157
rect 201 150 210 152
rect 225 157 234 159
rect 225 152 227 157
rect 232 152 234 157
rect 225 150 234 152
rect 249 157 258 159
rect 249 152 251 157
rect 256 152 258 157
rect 249 150 258 152
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
rect 131 5 136 10
rect 155 5 160 10
rect 179 5 184 10
rect 203 5 208 10
rect 227 5 232 10
rect 251 5 256 10
<< nsubdiffcont >>
rect 11 152 16 157
rect 35 152 40 157
rect 59 152 64 157
rect 83 152 88 157
rect 107 152 112 157
rect 131 152 136 157
rect 155 152 160 157
rect 179 152 184 157
rect 203 152 208 157
rect 227 152 232 157
rect 251 152 256 157
<< polysilicon >>
rect 19 143 25 148
rect 36 143 42 148
rect 53 143 59 148
rect 70 143 76 148
rect 87 143 93 148
rect 104 143 110 148
rect 121 143 127 148
rect 138 143 144 148
rect 155 143 161 148
rect 172 143 178 148
rect 189 143 195 148
rect 206 143 212 148
rect 223 143 229 148
rect 255 143 261 148
rect 19 78 25 109
rect 36 91 42 109
rect 30 89 42 91
rect 30 83 32 89
rect 38 83 42 89
rect 30 81 42 83
rect 12 76 25 78
rect 12 70 14 76
rect 20 70 25 76
rect 12 68 25 70
rect 19 36 25 68
rect 36 36 42 81
rect 53 65 59 109
rect 47 63 59 65
rect 47 57 49 63
rect 55 57 59 63
rect 47 55 59 57
rect 53 36 59 55
rect 70 91 76 109
rect 87 107 93 109
rect 104 107 110 109
rect 87 102 110 107
rect 70 89 82 91
rect 70 83 74 89
rect 80 83 82 89
rect 70 81 82 83
rect 70 36 76 81
rect 87 78 93 102
rect 121 91 127 109
rect 115 89 127 91
rect 115 83 117 89
rect 123 83 127 89
rect 115 81 127 83
rect 87 76 102 78
rect 87 70 94 76
rect 100 70 102 76
rect 87 68 102 70
rect 87 43 93 68
rect 87 38 110 43
rect 87 36 93 38
rect 104 36 110 38
rect 121 36 127 81
rect 138 52 144 109
rect 155 65 161 109
rect 149 63 161 65
rect 149 57 151 63
rect 157 57 161 63
rect 149 55 161 57
rect 133 50 144 52
rect 133 44 135 50
rect 141 44 144 50
rect 133 42 144 44
rect 138 36 144 42
rect 155 36 161 55
rect 172 78 178 109
rect 189 91 195 109
rect 189 89 201 91
rect 189 83 193 89
rect 199 83 201 89
rect 189 81 201 83
rect 172 76 184 78
rect 172 70 176 76
rect 182 70 184 76
rect 172 68 184 70
rect 172 36 178 68
rect 189 36 195 81
rect 206 52 212 109
rect 223 65 229 109
rect 255 65 261 109
rect 217 63 229 65
rect 217 57 219 63
rect 225 57 229 63
rect 217 55 229 57
rect 249 63 261 65
rect 249 57 251 63
rect 257 57 261 63
rect 249 55 261 57
rect 201 50 212 52
rect 201 44 203 50
rect 209 44 212 50
rect 201 42 212 44
rect 206 36 212 42
rect 223 36 229 55
rect 255 36 261 55
rect 19 14 25 19
rect 36 14 42 19
rect 53 14 59 19
rect 70 14 76 19
rect 87 14 93 19
rect 104 14 110 19
rect 121 14 127 19
rect 138 14 144 19
rect 155 14 161 19
rect 172 14 178 19
rect 189 14 195 19
rect 206 14 212 19
rect 223 14 229 19
rect 255 14 261 19
<< polycontact >>
rect 32 83 38 89
rect 14 70 20 76
rect 49 57 55 63
rect 74 83 80 89
rect 117 83 123 89
rect 94 70 100 76
rect 151 57 157 63
rect 135 44 141 50
rect 193 83 199 89
rect 176 70 182 76
rect 219 57 225 63
rect 251 57 257 63
rect 203 44 209 50
<< metal1 >>
rect 0 157 280 162
rect 0 151 11 157
rect 17 151 35 157
rect 41 151 59 157
rect 65 151 83 157
rect 89 151 107 157
rect 113 151 131 157
rect 137 151 155 157
rect 161 151 179 157
rect 185 151 203 157
rect 209 151 227 157
rect 233 151 251 157
rect 257 151 280 157
rect 0 150 280 151
rect 11 141 16 143
rect 11 104 16 111
rect 28 141 33 150
rect 28 109 33 111
rect 45 141 50 143
rect 45 104 50 111
rect 11 99 50 104
rect 62 141 67 143
rect 30 83 32 89
rect 38 83 40 89
rect 12 70 14 76
rect 20 70 22 76
rect 62 63 67 111
rect 96 141 101 150
rect 96 109 101 111
rect 113 141 118 143
rect 113 104 118 111
rect 130 141 135 150
rect 130 109 135 111
rect 147 141 152 143
rect 147 104 152 111
rect 113 99 152 104
rect 164 141 169 143
rect 72 83 74 89
rect 80 83 117 89
rect 123 83 125 89
rect 92 70 94 76
rect 100 70 102 76
rect 164 63 169 111
rect 215 141 220 150
rect 215 109 220 111
rect 232 141 237 143
rect 232 89 237 111
rect 247 141 252 150
rect 247 109 252 111
rect 264 141 269 143
rect 191 83 193 89
rect 199 83 201 89
rect 238 83 240 89
rect 174 70 176 76
rect 182 70 184 76
rect 47 57 49 63
rect 55 57 57 63
rect 62 57 151 63
rect 157 57 159 63
rect 164 57 219 63
rect 225 57 227 63
rect 11 41 50 46
rect 11 34 16 41
rect 11 19 16 21
rect 28 34 33 36
rect 28 12 33 21
rect 45 34 50 41
rect 45 19 50 21
rect 62 34 67 57
rect 133 44 135 50
rect 141 44 143 50
rect 62 19 67 21
rect 96 34 101 36
rect 96 12 101 21
rect 113 34 152 39
rect 113 33 118 34
rect 147 33 152 34
rect 113 19 118 21
rect 130 27 135 29
rect 130 12 135 21
rect 147 19 152 21
rect 164 34 169 57
rect 201 44 203 50
rect 209 44 211 50
rect 164 19 169 21
rect 215 34 220 36
rect 215 12 220 21
rect 232 34 237 83
rect 264 64 269 111
rect 264 63 272 64
rect 249 57 251 63
rect 257 57 259 63
rect 264 57 267 63
rect 273 57 275 63
rect 264 56 272 57
rect 232 19 237 21
rect 247 34 252 36
rect 247 12 252 21
rect 264 34 269 56
rect 264 19 269 21
rect 0 11 282 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 131 11
rect 137 5 155 11
rect 161 5 179 11
rect 185 5 203 11
rect 209 5 227 11
rect 233 5 251 11
rect 257 5 282 11
rect 0 0 282 5
<< via1 >>
rect 11 152 16 157
rect 16 152 17 157
rect 11 151 17 152
rect 35 152 40 157
rect 40 152 41 157
rect 35 151 41 152
rect 59 152 64 157
rect 64 152 65 157
rect 59 151 65 152
rect 83 152 88 157
rect 88 152 89 157
rect 83 151 89 152
rect 107 152 112 157
rect 112 152 113 157
rect 107 151 113 152
rect 131 152 136 157
rect 136 152 137 157
rect 131 151 137 152
rect 155 152 160 157
rect 160 152 161 157
rect 155 151 161 152
rect 179 152 184 157
rect 184 152 185 157
rect 179 151 185 152
rect 203 152 208 157
rect 208 152 209 157
rect 203 151 209 152
rect 227 152 232 157
rect 232 152 233 157
rect 227 151 233 152
rect 251 152 256 157
rect 256 152 257 157
rect 251 151 257 152
rect 32 83 38 89
rect 14 70 20 76
rect 74 83 80 89
rect 117 83 123 89
rect 94 70 100 76
rect 193 83 199 89
rect 232 83 238 89
rect 176 70 182 76
rect 49 57 55 63
rect 151 57 157 63
rect 135 44 141 50
rect 203 44 209 50
rect 251 57 257 63
rect 267 57 273 63
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 131 10 137 11
rect 131 5 136 10
rect 136 5 137 10
rect 155 10 161 11
rect 155 5 160 10
rect 160 5 161 10
rect 179 10 185 11
rect 179 5 184 10
rect 184 5 185 10
rect 203 10 209 11
rect 203 5 208 10
rect 208 5 209 10
rect 227 10 233 11
rect 227 5 232 10
rect 232 5 233 10
rect 251 10 257 11
rect 251 5 256 10
rect 256 5 257 10
<< metal2 >>
rect 10 157 18 158
rect 34 157 42 158
rect 58 157 66 158
rect 82 157 90 158
rect 106 157 114 158
rect 130 157 138 158
rect 154 157 162 158
rect 178 157 186 158
rect 202 157 210 158
rect 226 157 234 158
rect 250 157 258 158
rect 9 151 11 157
rect 17 151 19 157
rect 33 151 35 157
rect 41 151 43 157
rect 57 151 59 157
rect 65 151 67 157
rect 81 151 83 157
rect 89 151 91 157
rect 105 151 107 157
rect 113 151 115 157
rect 129 151 131 157
rect 137 151 139 157
rect 153 151 155 157
rect 161 151 163 157
rect 177 151 179 157
rect 185 151 187 157
rect 201 151 203 157
rect 209 151 211 157
rect 225 151 227 157
rect 233 151 235 157
rect 249 151 251 157
rect 257 151 259 157
rect 10 150 18 151
rect 34 150 42 151
rect 58 150 66 151
rect 82 150 90 151
rect 106 150 114 151
rect 130 150 138 151
rect 154 150 162 151
rect 178 150 186 151
rect 202 150 210 151
rect 226 150 234 151
rect 250 150 258 151
rect 31 89 39 90
rect 73 89 81 90
rect 116 89 124 90
rect 192 89 200 90
rect 231 89 239 90
rect 30 83 32 89
rect 38 83 74 89
rect 80 83 82 89
rect 115 83 117 89
rect 123 83 193 89
rect 199 83 201 89
rect 230 83 232 89
rect 238 83 240 89
rect 31 82 39 83
rect 73 82 81 83
rect 116 82 124 83
rect 192 82 200 83
rect 231 82 239 83
rect 13 76 21 77
rect 93 76 101 77
rect 175 76 183 77
rect 12 70 14 76
rect 20 70 94 76
rect 100 70 176 76
rect 182 70 184 76
rect 13 69 21 70
rect 93 69 101 70
rect 175 69 183 70
rect 48 63 56 64
rect 150 63 158 64
rect 250 63 258 64
rect 266 63 274 64
rect 47 57 49 63
rect 55 57 57 63
rect 149 57 151 63
rect 157 57 251 63
rect 257 57 259 63
rect 265 57 267 63
rect 273 57 275 63
rect 48 56 56 57
rect 150 56 158 57
rect 250 56 258 57
rect 266 56 274 57
rect 49 50 55 56
rect 251 55 257 56
rect 134 50 142 51
rect 202 50 210 51
rect 49 44 135 50
rect 141 44 203 50
rect 209 44 211 50
rect 134 43 142 44
rect 202 43 210 44
rect 135 42 141 43
rect 203 42 209 43
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 129 5 131 11
rect 137 5 139 11
rect 153 5 155 11
rect 161 5 163 11
rect 177 5 179 11
rect 185 5 187 11
rect 201 5 203 11
rect 209 5 211 11
rect 225 5 227 11
rect 233 5 235 11
rect 249 5 251 11
rect 257 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< labels >>
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 14 154 14 154 1 VDD
rlabel metal2 17 73 17 73 1 A
port 1 n
rlabel metal2 35 86 35 86 1 B
port 2 n
rlabel metal2 52 60 52 60 1 CI
port 3 n
rlabel metal2 270 60 270 60 1 CO
port 5 n
rlabel metal2 235 86 235 86 1 S
port 6 n
<< end >>
