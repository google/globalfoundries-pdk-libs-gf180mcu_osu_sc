magic
tech gf180mcuC
timestamp 1661875399
<< nwell >>
rect 0 61 80 123
<< nmos >>
rect 18 19 24 36
rect 35 19 41 36
rect 54 19 60 36
<< pmos >>
rect 21 70 27 104
rect 33 70 39 104
rect 52 70 58 104
<< ndiff >>
rect 8 28 18 36
rect 8 21 10 28
rect 15 21 18 28
rect 8 19 18 21
rect 24 26 35 36
rect 24 21 27 26
rect 32 21 35 26
rect 24 19 35 21
rect 41 28 54 36
rect 41 21 44 28
rect 51 21 54 28
rect 41 19 54 21
rect 60 32 70 36
rect 60 21 63 32
rect 68 21 70 32
rect 60 19 70 21
<< pdiff >>
rect 11 102 21 104
rect 11 72 13 102
rect 18 72 21 102
rect 11 70 21 72
rect 27 70 33 104
rect 39 102 52 104
rect 39 80 42 102
rect 49 80 52 102
rect 39 70 52 80
rect 58 102 68 104
rect 58 91 61 102
rect 66 91 68 102
rect 58 77 68 91
rect 58 70 69 77
<< ndiffc >>
rect 10 21 15 28
rect 27 21 32 26
rect 44 21 51 28
rect 63 21 68 32
<< pdiffc >>
rect 13 72 18 102
rect 42 80 49 102
rect 61 91 66 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
<< polysilicon >>
rect 21 104 27 109
rect 33 104 39 109
rect 52 104 58 109
rect 21 68 27 70
rect 16 64 27 68
rect 33 65 39 70
rect 16 52 22 64
rect 32 63 43 65
rect 32 57 35 63
rect 41 57 43 63
rect 32 55 43 57
rect 11 50 22 52
rect 11 44 14 50
rect 20 45 22 50
rect 33 45 39 55
rect 52 52 58 70
rect 47 50 60 52
rect 20 44 24 45
rect 11 42 24 44
rect 33 42 41 45
rect 47 44 49 50
rect 55 44 60 50
rect 47 42 60 44
rect 18 36 24 42
rect 35 36 41 42
rect 54 36 60 42
rect 18 14 24 19
rect 35 14 41 19
rect 54 14 60 19
<< polycontact >>
rect 35 57 41 63
rect 14 44 20 50
rect 49 44 55 50
<< metal1 >>
rect 0 118 80 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 80 118
rect 0 111 80 112
rect 13 102 18 111
rect 13 70 18 72
rect 42 102 49 104
rect 61 102 66 111
rect 61 89 66 91
rect 42 76 49 80
rect 42 70 62 76
rect 68 70 70 76
rect 62 69 69 70
rect 33 57 35 63
rect 41 57 43 63
rect 12 44 14 50
rect 20 44 22 50
rect 47 44 49 50
rect 55 44 57 50
rect 10 33 51 38
rect 10 28 15 33
rect 44 28 51 33
rect 10 19 15 21
rect 27 26 32 28
rect 27 12 32 21
rect 44 19 51 21
rect 63 32 68 69
rect 63 19 68 21
rect 0 11 80 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 80 11
rect 0 0 80 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 62 70 68 76
rect 35 57 41 63
rect 14 44 20 50
rect 49 44 55 50
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 61 76 69 77
rect 60 70 62 76
rect 68 70 70 76
rect 61 69 69 70
rect 33 63 43 64
rect 33 57 35 63
rect 41 57 43 63
rect 33 56 43 57
rect 12 50 22 51
rect 12 44 14 50
rect 20 44 22 50
rect 12 43 22 44
rect 47 50 57 51
rect 47 44 49 50
rect 55 44 57 50
rect 47 43 57 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 17 47 17 47 1 A0
port 5 n
rlabel metal2 38 60 38 60 1 A1
port 6 n
rlabel metal2 52 47 52 47 1 B
port 7 n
rlabel metal2 65 73 65 73 1 Y
port 4 n
<< end >>
