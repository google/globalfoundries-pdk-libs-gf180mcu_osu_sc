* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__nfet_01v8_lvt.0 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.417908+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.47213
+ k2 = -0.033282
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 161140.0
+ ua = -1.3015602e-9
+ ub = 2.67551e-18
+ uc = 7.0152e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03198837
+ a0 = 1.9598449
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.5317926
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11559919+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.1019079+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0047977
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.4345657e-5
+ alpha1 = 0.0
+ beta0 = 17.822982
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25364
+ kt2 = -0.034423
+ at = 333080.0
+ ute = -1.0777
+ ua1 = 2.6823e-9
+ ub1 = -2.4433e-18
+ uc1 = -1.9223e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.1 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.065634200e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(1))} lvth0 = 9.048380250e-08 wvth0 = 7.882214154e-08 pvth0 = -6.286814598e-13
+ k1 = 5.488515703e-01 lk1 = -6.119274088e-07 wk1 = -5.330614706e-07 pk1 = 4.251671636e-12
+ k2 = -5.971089207e-02 lk2 = 2.107955217e-07 wk2 = 1.836279421e-07 pk2 = -1.464607285e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.374663231e+04 lvsat = 6.970451310e-01 wvsat = 6.072091187e-01 pvsat = -4.843069571e-6
+ ua = -1.339853632e-09 lua = 3.054264999e-16 wua = 2.660627664e-16 pua = -2.122103322e-21
+ ub = 2.691095738e-18 lub = -1.243110679e-25 wub = -1.082897084e-25 pub = 8.637132995e-31
+ uc = 6.984327633e-11 luc = 2.462364538e-18 wuc = 2.145012044e-18 puc = -1.710850881e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.155047379e-02 lu0 = 3.492638310e-09 wu0 = 3.042502896e-09 pu0 = -2.426685098e-14
+ a0 = 1.997305793e+00 la0 = -2.987862100e-07 wa0 = -2.602782850e-07 pa0 = 2.075966587e-12
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.149843589e-01 lags = 1.340616906e-07 wags = 1.167836592e-07 pags = -9.314606265e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.120694636e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.815292095e-08 wvoff = -2.452453874e-08 pvoff = 1.956064948e-13
+ nfactor = {1.187777049e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -6.848880369e-07 wnfactor = -5.966188454e-07 pnfactor = 4.758602080e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.405322955e-01 lpclm = -1.120878562e-06 wpclm = -9.764183890e-07 ppclm = 7.787864250e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.886283880e-03 lpdiblc2 = 1.524535941e-08 wpdiblc2 = 1.328051920e-08 ppdiblc2 = -1.059247572e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.383516913e-04 lalpha0 = -4.307494292e-10 walpha0 = -3.752339263e-10 palpha0 = 2.992847034e-15
+ alpha1 = 0.0
+ beta0 = 1.812382841e+01 lbeta0 = -2.399535901e-06 wbeta0 = -2.090280837e-06 pbeta0 = 1.667197544e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.532233833e-01 lkt1 = -3.322914083e-09 wkt1 = -2.894652931e-09 pkt1 = 2.308760705e-14
+ kt2 = -3.413777779e-02 lkt2 = -2.274918103e-09 wkt2 = -1.981723930e-09 pkt2 = 1.580613098e-14
+ at = 6.161496924e+05 lat = -2.257749713e+00 wat = -1.966768223e+00 pat = 1.568684501e-5
+ ute = -9.503648401e-01 lute = -1.015618868e-06 wute = -8.847246908e-07 pute = 7.056519897e-12
+ ua1 = 2.422715740e-09 lua1 = 2.070431082e-15 wua1 = 1.803591442e-15 pua1 = -1.438535516e-20
+ ub1 = -1.556867822e-18 lub1 = -7.070138733e-24 wub1 = -6.158930775e-24 pub1 = 4.912332392e-29
+ uc1 = -1.093873687e-11 luc1 = -6.607486849e-17 wuc1 = -5.755906021e-17 puc1 = 4.590881863e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.2 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.272748110e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 8.136347530e-09 wvth0 = -1.576442831e-07 pvth0 = 3.114972211e-13
+ k1 = 3.599249359e-01 lk1 = 1.392354435e-07 wk1 = 1.066122941e-06 pk1 = -2.106605626e-12
+ k2 = 4.780166941e-03 lk2 = -4.561770435e-08 wk2 = -3.672558843e-07 pk2 = 7.256792645e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.501850562e+05 lvsat = -7.996552203e-01 wvsat = -1.214418237e+00 pvsat = 2.399629716e-6
+ ua = -1.300809062e-09 lua = 1.501872405e-16 wua = -5.321255328e-16 pua = 1.051453447e-21
+ ub = 2.626614252e-18 lub = 1.320640957e-25 wub = 2.165794168e-25 pub = -4.279500985e-31
+ uc = 6.801003316e-11 luc = 9.751247726e-18 wuc = -4.290024088e-18 puc = 8.476873096e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.075352180e-02 lu0 = 6.661279571e-09 wu0 = -6.085005793e-09 pu0 = 1.202366720e-14
+ a0 = 1.873713451e+00 la0 = 1.926107635e-07 wa0 = 5.205565699e-07 pa0 = -1.028593754e-12
+ keta = 1.823110268e-01 lketa = -7.248595268e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.674985624e-01 lags = 3.642769662e-06 wags = -2.335673184e-07 pags = 4.615173427e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.223648486e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.278101484e-08 wvoff = 4.904907748e-08 pvoff = -9.691852464e-14
+ nfactor = {6.880557574e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.301978831e-06 wnfactor = 1.193237691e-06 pnfactor = -2.357778015e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 8.336952366e-01 ldsub = -1.088198576e-6
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.108026385e-01 lpclm = 6.736065685e-07 wpclm = 1.952836778e-06 ppclm = -3.858707832e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 4.773555186e-03 lpdiblc2 = 7.741663056e-09 wpdiblc2 = -2.656103841e-08 ppdiblc2 = 5.248328385e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.460214106e-05 lalpha0 = 3.761848605e-10 walpha0 = 7.504678525e-10 palpha0 = -1.482886953e-15
+ alpha1 = 0.0
+ beta0 = 1.378943650e+01 lbeta0 = 1.483378959e-05 wbeta0 = 4.180561674e-06 pbeta0 = -8.260580840e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.544831132e-01 lkt1 = 1.685708985e-09 wkt1 = 5.789305862e-09 pkt1 = -1.143937892e-14
+ kt2 = -3.970410922e-02 lkt2 = 1.985653737e-08 wkt2 = 3.963447860e-09 pkt2 = -7.831574798e-15
+ at = 4.525514858e+04 lat = 1.209844826e-02 wat = 3.933536446e+00 pat = -7.772471341e-6
+ ute = -1.241970607e+00 lute = 1.437910814e-07 wute = 1.769449382e-06 pute = -3.496343505e-12
+ ua1 = 2.638520366e-09 lua1 = 1.212402678e-15 wua1 = -3.607182884e-15 pua1 = 7.127613019e-21
+ ub1 = -2.908579444e-18 lub1 = -1.695800907e-24 wub1 = 1.231786155e-23 pub1 = -2.433947853e-29
+ uc1 = -2.045321438e-11 luc1 = -2.824578165e-17 wuc1 = 1.151181204e-16 puc1 = -2.274676500e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.3 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.281499842e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 6.407049093e-9
+ k1 = 4.290139105e-01 lk1 = 2.719084048e-9
+ k2 = -1.426108485e-02 lk2 = -7.993142886e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.918426775e+04 lvsat = 5.198078759e-2
+ ua = -9.501342298e-10 lua = -5.427286938e-16
+ ub = 2.617706520e-18 lub = 1.496653283e-25
+ uc = 5.966524835e-11 luc = 2.624012527e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.824115950e-02 lu0 = -8.133918159e-9
+ a0 = 2.190574410e+00 la0 = -4.334906492e-07 wa0 = 3.388131789e-21
+ keta = -1.449161895e-01 lketa = -7.827490886e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 8.170574498e-01 lags = 1.302146209e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.170681977e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.315097581e-9
+ nfactor = {9.331405229e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.177035890e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.487975000e-05 lcit = -9.642142013e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.912122870e-04 leta0 = -1.802309185e-10
+ etab = -5.415949890e-04 letab = 8.218961851e-11
+ dsub = -5.153016090e-02 ldsub = 6.609625483e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.292314045e-01 lpclm = 1.716301278e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 7.015305875e-03 lpdiblc2 = 3.312075781e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.865945616e-04 lalpha0 = -1.201672640e-10
+ alpha1 = 0.0
+ beta0 = 2.119695075e+01 lbeta0 = 1.969118242e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.506826310e-01 lkt1 = -5.823853776e-9
+ kt2 = -4.595043715e-02 lkt2 = 3.219896904e-8
+ at = 3.099626020e+04 lat = 4.027329876e-2
+ ute = -1.324376050e+00 lute = 3.066201160e-7
+ ua1 = 3.273961280e-09 lua1 = -4.319679622e-17
+ ub1 = -3.908312750e-18 lub1 = 2.796221184e-25
+ uc1 = 1.127389820e-11 luc1 = -9.093696975e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.4 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.415412995e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -6.662205081e-9
+ k1 = 4.337989900e-01 lk1 = -1.950914290e-9
+ k2 = -1.718793358e-02 lk2 = -5.136684864e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.761046784e+04 lvsat = 5.351673761e-2
+ ua = -1.221602632e-09 lua = -2.777891065e-16
+ ub = 2.751298556e-18 lub = 1.928618127e-26
+ uc = 1.074233594e-10 luc = -2.036940321e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.407221921e-02 lu0 = -4.065240878e-9
+ a0 = 2.020645123e+00 la0 = -2.676481611e-7
+ keta = -4.305008473e-01 lketa = 2.004414379e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.933555805e+00 lags = -7.634503603e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.149696165e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.669872657e-10
+ nfactor = {1.346903917e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 4.138912047e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 7.840064260e-04 leta0 = -3.683883585e-10
+ etab = -8.332985405e-04 letab = 3.668776996e-10
+ dsub = 2.694433755e-01 ldsub = 3.477084254e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.127243800e-02 lpclm = 2.657145264e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.030333910e-02 lpdiblc2 = 1.031197554e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.816033686e-05 lalpha0 = 8.942277909e-11
+ alpha1 = 0.0
+ beta0 = 1.856086122e+01 lbeta0 = 2.769603395e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.506815870e-01 lkt1 = -5.824872667e-9
+ kt2 = -1.336252900e-03 lkt2 = -1.134224408e-8
+ at = 7.236385330e+04 lat = -9.940372813e-5
+ ute = -1.005059740e+00 lute = -5.016636747e-9
+ ua1 = 4.029867140e-09 lua1 = -7.809231203e-16
+ ub1 = -4.686309770e-18 lub1 = 1.038908310e-24
+ uc1 = -1.680361004e-10 luc1 = 8.406062335e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.5 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955659379e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.237523171e-8
+ k1 = 2.939492400e-01 lk1 = 6.461057422e-8
+ k2 = 1.411904655e-02 lk2 = -2.003724206e-08 pk2 = 1.262177448e-29
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.862158910e+04 lvsat = 1.495949445e-2
+ ua = -1.685639191e-09 lua = -5.693090631e-17
+ ub = 2.816927564e-18 lub = -1.194994509e-26
+ uc = 7.395486363e-11 luc = -4.440072643e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.785579897e-02 lu0 = -1.106535664e-9
+ a0 = 1.318301380e+00 la0 = 6.663234319e-8
+ keta = -1.362724654e-02 lketa = 2.030447647e-9
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.531102100e+00 lags = -5.719025195e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.186422400e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.014972382e-9
+ nfactor = {1.984499198e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.104277305e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -5.197693883e-03 leta0 = 2.478601904e-09 weta0 = -1.654361225e-24 peta0 = 6.779273404e-31
+ etab = 2.455547952e-02 letab = -1.171691122e-08 wetab = 7.031035207e-24 petab = 1.627025617e-30
+ dsub = 1.659631037e+00 ldsub = -3.139513920e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.407131060e-01 lpclm = -5.887649330e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 7.428100200e-03 lpdiblc2 = 1.471589710e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.283466402e-03 lalpha0 = 1.162835701e-09 walpha0 = -4.135903063e-25 palpha0 = 1.972152263e-31
+ alpha1 = 0.0
+ beta0 = 1.815423470e+01 lbeta0 = 2.963137290e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.539452660e-01 lkt1 = -4.271524647e-9
+ kt2 = -2.835108740e-02 lkt2 = 1.515466398e-9
+ at = 8.746446820e+04 lat = -7.286541390e-3
+ ute = -4.267743000e-01 lute = -2.802515919e-7
+ ua1 = 4.105298706e-09 lua1 = -8.168247741e-16
+ ub1 = -4.131849346e-18 lub1 = 7.750128712e-25
+ uc1 = 4.935840992e-11 luc1 = -1.940829382e-17 wuc1 = 2.465190329e-32
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.6 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.085981921e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.791486956e-8
+ k1 = 3.156315857e-01 lk1 = 5.971144821e-8
+ k2 = -4.315366053e-03 lk2 = -1.587198653e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.521236440e+05 lvsat = 2.870705142e-3
+ ua = -9.341333047e-10 lua = -2.267336613e-16
+ ub = 2.603968464e-18 lub = 3.616816349e-26
+ uc = 8.319096704e-11 luc = -6.526970211e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.935215995e-02 lu0 = -3.704138428e-9
+ a0 = 5.207179143e+00 la0 = -8.120595873e-7
+ keta = 2.463675731e-01 lketa = -5.671538185e-08 wketa = -6.617444900e-23 pketa = -1.577721810e-29
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.681894429e+00 lags = 6.059740461e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.639417362e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.225039357e-8
+ nfactor = {1.251539366e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.760400046e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.539000915e-01 leta0 = 3.607790865e-08 weta0 = 5.293955920e-23 peta0 = -2.208810535e-29
+ etab = -5.508974867e-02 letab = 6.278928090e-9
+ dsub = 1.548726549e-01 ldsub = 2.604876439e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.965795643e-01 lpclm = -1.166895196e-7
+ pdiblc1 = -9.689928571e-01 lpdiblc1 = 3.070644361e-07 ppdiblc1 = 2.019483917e-28
+ pdiblc2 = 1.446009071e-02 lpdiblc2 = -1.172885469e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.807445428e-03 lalpha0 = -1.117205827e-9
+ alpha1 = 0.0
+ beta0 = 3.632420408e+01 lbeta0 = -1.142367291e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.821762143e-01 lkt1 = -2.048774188e-8
+ kt2 = -3.510916857e-02 lkt2 = 3.042454839e-9
+ at = 1.366878571e+02 lat = 1.244517058e-2
+ ute = -1.139543429e+00 lute = -1.192014073e-7
+ ua1 = 1.541707280e-09 lua1 = -2.375812914e-16
+ ub1 = -1.995903100e-18 lub1 = 2.923958169e-25 pub1 = 3.503246161e-46
+ uc1 = -1.221356132e-10 luc1 = 1.934078071e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.7 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.499593467e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(1))} lvth0 = -1.985141613e-9
+ k1 = 1.011211867e+00 lk1 = -4.876429661e-8
+ k2 = -2.173785925e-01 lk2 = 1.735522364e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.819855190e+05 lvsat = -1.786254255e-3
+ ua = -3.496851673e-09 lua = 1.729222682e-16
+ ub = 4.579415850e-18 lub = -2.719028563e-25
+ uc = 1.863698448e-10 luc = -2.261771620e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.421071555e-02 lu0 = 2.166698265e-10
+ a0 = 0.0
+ keta = 1.569286063e-01 lketa = -4.276737498e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.005218833e+00 lags = 3.096873294e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.193483187e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 5.296050099e-9
+ nfactor = {7.234594002e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.583940752e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 6.763735176e-02 leta0 = 1.529144370e-9
+ etab = -7.707727382e-02 letab = 9.707882638e-9
+ dsub = 5.818051642e-01 ldsub = -4.053136044e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.682441667e-02 lpclm = 9.591795721e-9
+ pdiblc1 = 3.583688214e+00 lpdiblc1 = -4.029261770e-7
+ pdiblc2 = 6.473580283e-02 lpdiblc2 = -7.957785852e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.687407636e-03 lalpha0 = -1.627859335e-10
+ alpha1 = 0.0
+ beta0 = 3.124083183e+01 lbeta0 = -3.496153888e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.951193167e-01 lkt1 = -2.874265066e-9
+ kt2 = 2.122778000e-02 lkt2 = -5.743292291e-9
+ at = 6.394335000e+04 lat = 2.494521618e-3
+ ute = -2.841387833e+00 lute = 1.462012276e-7
+ ua1 = -2.429022070e-09 lua1 = 3.816539507e-16 wua1 = 9.860761315e-32 pua1 = 1.293043786e-37
+ ub1 = 2.444379600e-18 lub1 = -4.000662701e-25 wub1 = 1.469367939e-39 pub1 = -8.758115402e-47
+ uc1 = 5.214877500e-12 luc1 = -5.195283211e-19
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.8 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.906886357e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 1.891201432e-7
+ k1 = 6.562101846e-01 wk1 = -1.278989123e-6
+ k2 = -9.669357138e-02 wk2 = 4.405835979e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.854532308e+04 wvsat = 1.456893625e+0
+ ua = -1.393438690e-09 wua = 6.383717507e-16
+ ub = 2.712905292e-18 wub = -2.598224910e-25
+ uc = 6.941127077e-11 wuc = 5.146586695e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.093771351e-02 wu0 = 7.299961309e-9
+ a0 = 2.049725856e+00 wa0 = -6.244928844e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.914641225e-01 wags = 2.802022619e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.071302200e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = -5.884240377e-8
+ nfactor = {1.307936122e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -1.431484089e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.371830215e-01 wpclm = -2.342747634e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.115864615e-04 wpdiblc2 = 3.186431687e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.139238281e-04 walpha0 = -9.003091326e-10
+ alpha1 = 0.0
+ beta0 = 1.854481110e+01 wbeta0 = -5.015268597e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526404000e-01 wkt1 = -6.945220800e-9
+ kt2 = -3.373865846e-02 wkt2 = -4.754805009e-9
+ at = 1.012256938e+06 wat = -4.718921368e+0
+ ute = -7.721812308e-01 wute = -2.122744409e-6
+ ua1 = 2.059472308e-09 wua1 = 4.327406806e-15
+ ub1 = -3.164587692e-19 wub1 = -1.477729287e-23
+ uc1 = 6.536615385e-13 wuc1 = -1.381030444e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.9 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.906886357e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 1.891201432e-7
+ k1 = 6.562101846e-01 wk1 = -1.278989123e-6
+ k2 = -9.669357138e-02 wk2 = 4.405835979e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.854532308e+04 wvsat = 1.456893625e+0
+ ua = -1.393438690e-09 wua = 6.383717507e-16
+ ub = 2.712905292e-18 wub = -2.598224910e-25
+ uc = 6.941127077e-11 wuc = 5.146586695e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.093771351e-02 wu0 = 7.299961309e-9
+ a0 = 2.049725856e+00 wa0 = -6.244928844e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.914641225e-01 wags = 2.802022619e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.071302200e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = -5.884240377e-8
+ nfactor = {1.307936122e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -1.431484089e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.371830215e-01 wpclm = -2.342747634e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.115864615e-04 wpdiblc2 = 3.186431687e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.139238281e-04 walpha0 = -9.003091326e-10
+ alpha1 = 0.0
+ beta0 = 1.854481110e+01 wbeta0 = -5.015268597e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.526404000e-01 wkt1 = -6.945220800e-9
+ kt2 = -3.373865846e-02 wkt2 = -4.754805009e-9
+ at = 1.012256938e+06 wat = -4.718921368e+0
+ ute = -7.721812308e-01 wute = -2.122744409e-6
+ ua1 = 2.059472308e-09 wua1 = 4.327406806e-15
+ ub1 = -3.164587692e-19 wub1 = -1.477729287e-23
+ uc1 = 6.536615385e-13 wuc1 = -1.381030444e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.10 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.387074751e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 2.066744953e-07 wvth0 = 4.577215666e-07 pvth0 = -1.067945829e-12
+ k1 = 1.043658291e+00 lk1 = -1.540474298e-06 wk1 = -3.684456410e-06 pk1 = 9.564017660e-12
+ k2 = -2.346599121e-01 lk2 = 5.485472722e-07 wk2 = 1.296373785e-06 pk2 = -3.402578993e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.335375596e+05 lvsat = 3.379248828e-01 wvsat = 2.841286497e+00 pvsat = -5.504276840e-6
+ ua = -1.628156003e-09 lua = 9.332242992e-16 wua = 1.742281014e-15 pua = -4.389088037e-21
+ ub = 2.607033192e-18 lub = 4.209421767e-25 wub = 3.526286227e-25 pub = -2.435075005e-30
+ uc = 1.251089846e-10 luc = -2.214513252e-16 wuc = -4.010135385e-16 puc = 1.614872350e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.453968505e-02 lu0 = 2.543824125e-08 wu0 = 3.708873192e-08 pu0 = -1.184386625e-13
+ a0 = 1.998634175e+00 la0 = 2.031379692e-07 wa0 = -3.473926242e-07 pa0 = -1.101736780e-12
+ keta = 1.026209329e-01 lketa = -4.080156980e-07 wketa = 5.536867724e-07 pketa = -2.201430923e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.735004679e-01 lags = 4.631840963e-06 wags = 1.892533921e-06 pags = -6.410550058e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.695778636e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -8.020458739e-08 wvoff = -1.969591909e-07 pvoff = 5.491454397e-13
+ nfactor = {1.764527776e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.815385585e-06 wnfactor = -6.286089894e-06 pnfactor = 1.930166995e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.661279615e-06 lcit = 5.034061469e-11 wcit = 8.797057077e-11 pcit = -3.497665908e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 1.184116408e+00 ldsub = -2.481455632e-06 wdsub = -2.434726299e-06 pdsub = 9.680350028e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.827566924e-01 lpclm = 6.139913634e-07 wpclm = -1.476413453e-06 ppclm = -3.444501387e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.933641797e-03 lpdiblc2 = 3.238502030e-08 wpdiblc2 = 6.172856623e-08 ppdiblc2 = -1.187387623e-13
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.094116620e-04 lalpha0 = -3.796548533e-10 walpha0 = -1.848180051e-09 palpha0 = 3.768687378e-15
+ alpha1 = 0.0
+ beta0 = 1.587877845e+01 lbeta0 = 1.060001253e-05 wbeta0 = -1.033618616e-05 pbeta0 = 2.115570220e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.794415474e-01 lkt1 = 1.065600221e-07 wkt1 = 1.792005069e-07 pkt1 = -7.401061062e-13
+ kt2 = -1.800388894e-02 lkt2 = -6.256065688e-08 wkt2 = -1.468096827e-07 pkt2 = 5.648030909e-13
+ at = 1.978932325e+06 lat = -3.843453004e+00 wat = -9.501652578e+00 pat = 1.901590015e-5
+ ute = -5.425074425e-01 lute = -9.131714985e-07 wute = -3.090420687e-06 pute = 3.847432499e-12
+ ua1 = -6.951433487e-10 lua1 = 1.095221412e-14 wua1 = 1.955511261e-14 pua1 = -6.054459688e-20
+ ub1 = 5.349391812e-18 lub1 = -2.252713862e-23 wub1 = -4.505852274e-23 pub1 = 1.203966559e-28
+ uc1 = 2.359887021e-11 luc1 = -9.122900240e-17 wuc1 = -1.909557633e-16 puc1 = 2.101397678e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.11 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.501238099e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.347861141e-08 wvth0 = -1.526741411e-07 pvth0 = 1.381655692e-13
+ k1 = 1.098075300e-01 lk1 = 3.047681127e-07 wk1 = 2.217845931e-06 pk1 = -2.098636651e-12
+ k2 = 1.011602926e-01 lk2 = -1.150166613e-07 wk2 = -8.019477308e-07 pk2 = 7.435994056e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.224886622e+03 lvsat = 5.978532721e-02 wvsat = 8.309378008e-02 pvsat = -5.422594129e-8
+ ua = -8.783334105e-10 lua = -5.483876523e-16 wua = -4.988720921e-16 pua = 3.931844360e-23
+ ub = 2.780493269e-18 lub = 7.819373686e-26 wub = -1.131042332e-24 pub = 4.965846175e-31
+ uc = -8.467754604e-11 luc = 1.930763700e-16 wuc = 1.002893735e-15 puc = -1.159178228e-21
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.324278166e-02 lu0 = -1.151814250e-08 wu0 = -3.475127073e-08 pu0 = 2.351359072e-14
+ a0 = 2.503276966e+00 la0 = -7.940109526e-07 wa0 = -2.172657356e-06 pa0 = 2.504895068e-12
+ keta = 1.545693683e-01 lketa = -5.106632091e-07 wketa = -2.080825656e-06 pketa = 3.004233910e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 8.744391799e-01 lags = 1.573189616e-06 wags = -3.986882604e-07 pags = -1.883209590e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.422342947e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.901902929e-08 wvoff = 1.748540418e-07 pvoff = -1.855389175e-13
+ nfactor = {-2.134306463e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.092961359e-06 wnfactor = 7.966376483e-06 pnfactor = -8.860490989e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.020230923e-05 lcit = -3.435569369e-11 wcit = -1.759411415e-10 pcit = 1.717097571e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 7.564320637e-04 leta0 = -5.066969362e-10 weta0 = -1.147947008e-09 peta0 = 2.268285891e-15
+ etab = -5.889721664e-04 letab = 1.758045523e-10 wetab = 3.291766289e-10 petab = -6.504365598e-16
+ dsub = 1.838639089e-01 ldsub = -5.050067068e-07 wdsub = -1.635517997e-06 pdsub = 8.101154384e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.250925600e+00 lpclm = -1.101466990e-06 wpclm = -7.098731270e-06 ppclm = 7.664917504e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.059719894e-02 lpdiblc2 = -4.230994463e-09 wpdiblc2 = -2.488699303e-08 ppdiblc2 = 5.240925206e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.606289833e-04 lalpha0 = -8.566771924e-11 walpha0 = 1.804088381e-10 palpha0 = -2.397028372e-16
+ alpha1 = 0.0
+ beta0 = 2.068289695e+01 lbeta0 = 1.107314584e-06 wbeta0 = 3.571645802e-06 pbeta0 = -6.325478373e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.145610854e-01 lkt1 = -2.164052685e-08 wkt1 = -2.509724988e-07 pkt1 = 1.098942445e-13
+ kt2 = -1.422016137e-01 lkt2 = 1.828478374e-07 wkt2 = 6.687531747e-07 pkt2 = -1.046708337e-12
+ at = 2.886737031e+01 lat = 6.676128345e-02 wat = 2.151614454e-01 pat = -1.840385176e-7
+ ute = -1.405967708e+00 lute = 7.929828131e-07 wute = 5.668988396e-07 pute = -3.379248019e-12
+ ua1 = 3.791858500e-09 lua1 = 2.086122817e-15 wua1 = -3.598349883e-15 pua1 = -1.479451267e-20
+ ub1 = -4.764213727e-18 lub1 = -2.543159755e-24 wub1 = 5.946799988e-24 pub1 = 1.961268845e-29
+ uc1 = 1.699225986e-10 luc1 = -3.803573735e-16 wuc1 = -1.102291170e-15 puc1 = 2.010892965e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.12 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.424712187e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -6.010065057e-09 wvth0 = -6.461078861e-09 pvth0 = -4.531068884e-15
+ k1 = 4.497027542e-01 lk1 = -2.695263127e-08 wk1 = -1.104993533e-07 pk1 = 1.737119296e-13
+ k2 = -1.909791244e-02 lk2 = 2.349333997e-09 wk2 = 1.327053315e-08 pk2 = -5.201285905e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.504710501e+05 lvsat = -8.001576602e-02 wvsat = -9.231153254e-01 pvsat = 9.277838352e-7
+ ua = -6.384869914e-10 lua = -7.824657650e-16 wua = -4.051487472e-15 pua = 3.506493423e-21
+ ub = 2.416060118e-18 lub = 4.338622712e-25 wub = 2.329236668e-24 pub = -2.880474673e-30
+ uc = 1.378981169e-10 luc = -2.414634830e-17 wuc = -2.117386152e-16 puc = 2.624221452e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.981974313e-02 lu0 = -8.177428043e-09 wu0 = -3.993379617e-08 pu0 = 2.857147642e-14
+ a0 = 2.170538518e+00 la0 = -4.692748649e-07 wa0 = -1.041459314e-06 pa0 = 1.400902338e-12
+ keta = -6.878723148e-01 lketa = 3.115177515e-07 wketa = 1.788216956e-06 pketa = -7.717582269e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.708129977e-01 lags = 1.967108588e-06 wags = 1.711113702e-05 pags = -1.897192358e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.108792756e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.581901611e-09 wvoff = -2.841968880e-08 pvoff = 1.284607991e-14
+ nfactor = {1.772922212e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.543802876e-07 wnfactor = -2.959975114e-06 pnfactor = 1.803081852e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.291689863e-04 leta0 = -1.873044940e-10 weta0 = 2.465410829e-09 peta0 = -1.258170690e-15
+ etab = -7.400703663e-04 letab = 3.232688405e-10 wetab = -6.477493539e-10 petab = 3.029943531e-16
+ dsub = -1.603029450e+00 ldsub = 1.238911867e-06 wdsub = 1.300994119e-05 pdsub = -6.192081509e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.762763149e-01 lpclm = 6.817907193e-07 wpclm = 3.717206937e-06 ppclm = -2.890897389e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 6.682104373e-04 lpdiblc2 = 5.459201868e-09 wpdiblc2 = 6.694487395e-08 ppdiblc2 = -3.721405852e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.076349711e-04 lalpha0 = 1.761444871e-10 walpha0 = 5.521897589e-10 palpha0 = -6.025424269e-16
+ alpha1 = 0.0
+ beta0 = 1.830440783e+01 lbeta0 = 3.428601033e-06 wbeta0 = 1.781838139e-06 pbeta0 = -4.578715585e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.182503416e-01 lkt1 = -1.803999725e-08 wkt1 = -2.253322930e-07 pkt1 = 8.487068561e-14
+ kt2 = 8.950120937e-02 lkt2 = -4.328253281e-08 wkt2 = -6.311386879e-07 pkt2 = 2.219211261e-13
+ at = 1.148750153e+04 lat = 5.557822944e-02 wat = 4.229688921e-01 pat = -3.868481952e-7
+ ute = -2.623470978e-01 lute = -3.231337214e-07 wute = -5.160367438e-06 pute = 2.210277504e-12
+ ua1 = 9.336718781e-09 lua1 = -3.325383575e-15 wua1 = -3.687200520e-14 pua1 = 1.767891124e-20
+ ub1 = -1.212596015e-17 lub1 = 4.641536672e-24 wub1 = 5.169069087e-23 pub1 = -2.503106186e-29
+ uc1 = -5.217161532e-10 luc1 = 2.946474663e-16 wuc1 = 2.457369007e-15 puc1 = -1.463157385e-21
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.13 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.046381253e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.559840423e-08 wvth0 = -6.303355817e-08 pvth0 = 2.239460264e-14
+ k1 = 2.736310936e-01 lk1 = 5.684867557e-08 wk1 = 1.411704813e-07 pk1 = 5.392967182e-14
+ k2 = 2.513163981e-02 lk2 = -1.870172140e-08 wk2 = -7.651549795e-08 pk2 = -9.279197553e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.952846699e+05 lvsat = 8.454666889e-02 wvsat = 2.042060687e+00 pvsat = -4.834916880e-7
+ ua = -2.029160092e-09 lua = -1.205749030e-16 wua = 2.386783217e-15 pua = 4.421984890e-22
+ ub = 3.206404926e-18 lub = 5.769765971e-26 wub = -2.706088712e-24 pub = -4.839115581e-31
+ uc = 1.347648575e-10 luc = -2.265507346e-17 wuc = -4.225078371e-16 puc = 1.265578257e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.660475222e-02 lu0 = -1.887753122e-09 wu0 = 8.692272785e-09 pu0 = 5.427898902e-15
+ a0 = 4.105362724e-01 la0 = 3.683982041e-07 wa0 = 6.307151968e-06 pa0 = -2.096669201e-12
+ keta = -1.305217443e-01 lketa = 4.624674752e-08 wketa = 8.121829703e-07 pketa = -3.072148516e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 8.764768139e+00 lags = -1.980399361e-06 wags = -4.331151164e-05 pags = 9.786236055e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.231742978e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.269914194e-09 wvoff = 3.148873777e-08 pvoff = -1.566733571e-14
+ nfactor = {2.098751310e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -6.980714917e-10 wnfactor = -7.938236699e-07 pnfactor = 7.721020721e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.021461833e-02 leta0 = 4.878606545e-09 weta0 = 3.485759816e-08 peta0 = -1.667523225e-14
+ etab = -4.249328683e-02 letab = 2.019571222e-08 wetab = 4.658548286e-07 petab = -2.217289076e-13
+ dsub = 1.820262607e+00 ldsub = -3.904039879e-07 wdsub = -1.116068150e-06 pdsub = 5.311926360e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.315063217e+00 lpclm = -2.183923309e-07 wpclm = -4.685384571e-06 ppclm = 1.108316040e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 1.276766690e-02 lpdiblc2 = -2.995344368e-10 wpdiblc2 = -3.709930945e-08 ppdiblc2 = 1.230577057e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.448795377e-03 lalpha0 = 2.242319782e-09 walpha0 = 1.504470572e-08 palpha0 = -7.500255397e-15
+ alpha1 = 0.0
+ beta0 = 1.851521036e+01 lbeta0 = 3.328269572e-06 wbeta0 = -2.508058894e-06 pbeta0 = -2.536939092e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.780772817e-01 lkt1 = -3.716036509e-08 wkt1 = -5.271307546e-07 pkt1 = 2.285116634e-13
+ kt2 = 6.870079521e-03 lkt2 = -3.954246557e-09 wkt2 = -2.447166678e-07 pkt2 = 3.800356561e-14
+ at = 1.790869369e+05 lat = -2.419072180e-02 wat = -6.365929122e-01 pat = 1.174502455e-7
+ ute = 1.632015465e+00 lute = -1.224755583e-06 wute = -1.430447129e-05 pute = 6.562413731e-12
+ ua1 = 8.772002011e-09 lua1 = -3.056606628e-15 wua1 = -3.242425456e-14 pua1 = 1.556200432e-20
+ ub1 = -7.742786767e-18 lub1 = 2.555365298e-24 wub1 = 2.508879320e-23 pub1 = -1.236988866e-29
+ uc1 = 3.030103002e-10 luc1 = -9.788108918e-17 wuc1 = -1.762373333e-15 puc1 = 5.452289821e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.14 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.118621589e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.982567463e-08 wvth0 = -2.267804122e-08 pvth0 = 1.327627359e-14
+ k1 = 1.682851083e-01 lk1 = 8.065160094e-08 wk1 = 1.023763325e-06 pk1 = -1.454921812e-13
+ k2 = 3.885495103e-02 lk2 = -2.180250357e-08 wk2 = -2.999473631e-07 pk2 = 4.120523238e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.900498318e+05 lvsat = -2.519661753e-03 wvsat = -2.635111525e-01 pvsat = 3.745226918e-8
+ ua = -3.170460283e-09 lua = 1.373018754e-16 wua = 1.553799985e-14 pua = -2.529318909e-21
+ ub = 4.758410537e-18 lub = -2.929780080e-25 wub = -1.496906352e-23 pub = 2.286907600e-30
+ uc = -1.275427629e-11 luc = 1.067687481e-17 wuc = 6.666275507e-16 puc = -1.195323152e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.105891285e-02 lu0 = -6.346707162e-10 wu0 = 1.271014808e-07 pu0 = -2.132666166e-14
+ a0 = 6.587983926e+00 la0 = -1.027396093e-06 wa0 = -9.593831633e-06 pa0 = 1.496158043e-12
+ keta = 6.886116130e-01 lketa = -1.388364346e-07 wketa = -3.072711589e-06 pketa = 5.705770742e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.749845442e+00 lags = 6.213275777e-07 wags = 4.721236442e-07 pags = -1.066763374e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.745077203e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.586870100e-08 wvoff = 7.341245702e-08 pvoff = -2.514000007e-14
+ nfactor = {2.563830907e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 4.155850276e-07 wnfactor = 6.914345801e-06 pnfactor = -9.695588197e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -2.241036374e-07 lcit = 1.180386217e-12 wcit = 3.629707207e-11 pcit = -8.201323435e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -5.857628930e-02 leta0 = 1.580592587e-08 weta0 = -6.623097778e-07 peta0 = 1.408497363e-13
+ etab = 1.720249857e-01 letab = -2.827469146e-08 wetab = -1.577993174e-06 petab = 2.400785486e-13
+ dsub = -4.412068082e-01 ldsub = 1.205750265e-07 wdsub = 4.141560110e-06 pdsub = -6.567684693e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 7.310477266e-01 lpclm = -8.643403085e-08 wpclm = 1.150115208e-06 ppclm = -2.102151355e-13
+ pdiblc1 = -9.690011940e-01 lpdiblc1 = 3.070663198e-07 wpdiblc1 = 5.792441349e-11 ppdiblc1 = -1.308802123e-17
+ pdiblc2 = -1.399733861e-02 lpdiblc2 = 5.748018559e-09 wpdiblc2 = 1.977222189e-07 ppdiblc2 = -4.075215377e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.098787927e-02 lalpha0 = -3.505096855e-09 walpha0 = -9.157765437e-08 palpha0 = 1.659106686e-14
+ alpha1 = 0.0
+ beta0 = 5.064741493e+01 lbeta0 = -3.932002052e-06 wbeta0 = -9.951766904e-05 pbeta0 = 1.938238232e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.809161004e-01 lkt1 = 8.671065990e-09 wkt1 = 1.380844729e-06 pkt1 = -2.025953971e-13
+ kt2 = -8.864338002e-02 lkt2 = 1.762701963e-08 wkt2 = 3.719557011e-07 pkt2 = -1.013335561e-13
+ at = 7.209416075e+04 lat = -1.570404195e-05 wat = -4.999605217e-01 pat = 8.657815686e-8
+ ute = -6.188275033e+00 lute = 5.422390548e-07 wute = 3.507858718e-05 pute = -4.595688331e-12
+ ua1 = -1.385078990e-08 lua1 = 2.055013205e-15 wua1 = 1.069470704e-13 pua1 = -1.592894656e-20
+ ub1 = 1.150465572e-17 lub1 = -1.793594333e-24 wub1 = -9.380188271e-23 pub1 = 1.449345956e-29
+ uc1 = -4.351785849e-10 luc1 = 6.891268941e-17 wuc1 = 2.175022567e-15 puc1 = -3.444256217e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.15 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.05e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.645687442e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.665266596e-09 wvth0 = -1.015060938e-07 pvth0 = 2.556950838e-14
+ k1 = 1.589330356e+00 lk1 = -1.409604054e-07 wk1 = -4.016767262e-06 pk1 = 6.405785639e-13
+ k2 = -3.863594104e-01 lk2 = 4.450967610e-08 wk2 = 1.174078723e-06 pk2 = -1.886691357e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.521302627e+05 lvsat = 3.393895041e-03 wvsat = 2.074343203e-01 pvsat = -3.599167731e-8
+ ua = -6.864350754e-09 lua = 7.133640943e-16 wua = 2.339738362e-14 pua = -3.754989808e-21
+ ub = 1.065127934e-17 lub = -1.211970898e-24 wub = -4.218730751e-23 pub = 6.531592751e-30
+ uc = 4.100475213e-10 luc = -5.525906552e-17 wuc = -1.554112496e-15 puc = 2.267920951e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.010834965e-02 lu0 = -4.864303858e-10 wu0 = -4.097676176e-08 pu0 = 4.885140275e-15
+ a0 = 0.0
+ keta = 5.960802604e-01 lketa = -1.244061701e-07 wketa = -3.051225693e-06 pketa = 5.672263486e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.171303655e+00 lags = 9.824375992e-09 wags = -1.153957340e-06 pags = 1.469109921e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-4.190333247e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 5.400246901e-08 wvoff = 2.082211422e-06 pvoff = -3.384121986e-13
+ nfactor = {-2.636019729e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.666552473e-07 wnfactor = 2.334166099e-05 pnfactor = -3.531398623e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.718957515e-05 lcit = -1.535276991e-12 wcit = -8.469316817e-11 pcit = 1.066710453e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.111874360e-01 leta0 = 5.520063420e-08 weta0 = 2.632074625e-06 peta0 = -3.729095113e-13
+ etab = -1.756825561e-01 letab = 2.595029969e-08 wetab = 6.851095014e-07 petab = -1.128523136e-13
+ dsub = 6.340608263e-01 ldsub = -4.711296107e-08 wdsub = -3.630723397e-07 pdsub = 4.572896119e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.369884534e+00 lpclm = -1.860606310e-07 wpclm = -8.914701697e-06 ppclm = 1.359393061e-12
+ pdiblc1 = 8.993563655e+00 lpdiblc1 = -1.246595668e-06 wpdiblc1 = -3.758781457e-05 ppdiblc1 = 5.861815627e-12
+ pdiblc2 = 1.271247206e-01 lpdiblc2 = -1.625996658e-08 wpdiblc2 = -4.334782007e-07 ppdiblc2 = 5.768355168e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.684812109e-03 lalpha0 = 8.104593659e-10 walpha0 = 5.817018278e-08 palpha0 = -6.762108340e-15
+ alpha1 = 0.0
+ beta0 = 2.028701882e+01 lbeta0 = 8.027017212e-07 wbeta0 = 7.610709275e-05 pbeta0 = -8.006299281e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 9.169068374e-02 lkt1 = -6.503196200e-08 wkt1 = -2.687555883e-06 pkt1 = 4.318716783e-13
+ kt2 = 3.628031166e-01 lkt2 = -5.277606152e-08 wkt2 = -2.373265438e-06 pkt2 = 3.267836806e-13
+ at = -7.713296612e+04 lat = 2.325626639e-02 wat = 9.801982444e-01 pat = -1.442526027e-7
+ ute = -4.278255164e+00 lute = 2.443714563e-07 wute = 9.983354214e-06 pute = -6.820867490e-13
+ ua1 = -6.873444496e-09 lua1 = 9.668961886e-16 wua1 = 3.087984701e-14 pua1 = -4.066263069e-21
+ ub1 = 5.970576591e-18 lub1 = -9.305546923e-25 wub1 = -2.450001669e-23 pub1 = 3.685833557e-30
+ uc1 = -2.592159638e-10 luc1 = 4.147131865e-17 wuc1 = 1.837265485e-15 puc1 = -2.917524047e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.16 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4285278+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.40031
+ k2 = -0.008541591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26571325e-9
+ ub = 2.66092e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03239829
+ a0 = 1.9247773
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.547527
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11890341+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.02152474+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.17 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4285278+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.40031
+ k2 = -0.008541591
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 242950.0
+ ua = -1.26571325e-9
+ ub = 2.66092e-18
+ uc = 7.0441e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03239829
+ a0 = 1.9247773
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.547527
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11890341+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.02152474+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.068446
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25403
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.18 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.302884208e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -7.000140464e-9
+ k1 = 3.064721345e-01 lk1 = 3.730946613e-7
+ k2 = 2.471859627e-02 lk2 = -1.322408416e-07 pk2 = 3.231174268e-27
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.349471337e+05 lvsat = -7.633710035e-01 pvsat = -5.421010862e-20
+ ua = -1.279560362e-09 lua = 5.505542420e-17
+ ub = 2.677587138e-18 lub = -6.626770832e-26
+ uc = 4.487418295e-11 luc = 1.016523862e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.196039972e-02 lu0 = 1.741029857e-9
+ a0 = 1.929127848e+00 la0 = -1.729756097e-8
+ keta = 2.134026000e-01 lketa = -8.484780675e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.948422205e-01 lags = 3.349217902e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.263653876e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.966844976e-8
+ nfactor = {5.068067088e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.046493156e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.493987500e-05 lcit = -1.964069601e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 6.969762922e-01 ldsub = -5.446108888e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.735584150e-02 lpclm = -7.518458431e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.417011710e-03 lpdiblc2 = 8.627764942e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.037226179e-05 lalpha0 = 3.743842380e-10
+ alpha1 = 0.0
+ beta0 = 1.381071399e+01 lbeta0 = 1.483284610e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.435871042e-01 lkt1 = -4.152043136e-8
+ kt2 = -4.737757495e-02 lkt2 = 5.044516362e-8
+ at = 7.784137337e+04 lat = -3.875109322e-2
+ ute = -1.160838912e+00 lute = -1.433770808e-7
+ ua1 = 3.217444208e-09 lua1 = -1.161550762e-15
+ ub1 = -3.665918860e-18 lub1 = 1.561828146e-24
+ uc1 = -1.460756502e-11 luc1 = -4.918423094e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.19 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.195767629e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.416556009e-8
+ k1 = 5.535542150e-01 lk1 = -1.151271756e-07 wk1 = -5.421010862e-20
+ k2 = -5.929343500e-02 lk2 = 3.376273163e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.385029280e+04 lvsat = 4.893579914e-2
+ ua = -9.781477547e-10 lua = -5.405208168e-16
+ ub = 2.554194283e-18 lub = 1.775504030e-25
+ uc = 1.159814647e-10 luc = -3.885204703e-17 wuc = 1.262177448e-29
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.628974630e-02 lu0 = -6.813542516e-9
+ a0 = 2.068571612e+00 la0 = -2.928314672e-07 wa0 = -2.168404345e-19
+ keta = -2.617622955e-01 lketa = 9.042400779e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 7.946696200e-01 lags = 1.196396981e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.072494924e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -8.103603264e-9
+ nfactor = {1.380482216e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.201540387e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.267507895e-04 leta0 = -5.285822251e-11
+ etab = -5.231104960e-04 letab = 4.566518457e-11
+ dsub = -1.433705843e-01 ldsub = 1.115872522e-06 pdsub = -5.169878828e-26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.693887798e-01 lpclm = 4.321299501e-07 ppclm = -6.462348536e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 5.617808580e-03 lpdiblc2 = 6.255050366e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.967251894e-04 lalpha0 = -1.336274706e-10
+ alpha1 = 0.0
+ beta0 = 2.139751195e+01 lbeta0 = -1.582873317e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.647756710e-01 lkt1 = 3.471171125e-10
+ kt2 = -8.397457100e-03 lkt2 = -2.657760024e-8
+ at = 4.307837625e+04 lat = 2.993885095e-2
+ ute = -1.292542570e+00 lute = 1.168627612e-7
+ ua1 = 3.071900540e-09 lua1 = -8.739637520e-16
+ ub1 = -3.574377795e-18 lub1 = 1.380947579e-24 wub1 = 3.761581923e-37
+ uc1 = -5.062385405e-11 luc1 = 2.198215536e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.20 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.411784859e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -6.916641465e-9
+ k1 = 4.275940400e-01 lk1 = 7.803657162e-9
+ k2 = -1.644274375e-02 lk2 = -8.057400507e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.422589378e+04 lvsat = 1.056152534e-1
+ ua = -1.449108734e-09 lua = -8.088644864e-17
+ ub = 2.882093865e-18 lub = -1.424631935e-25
+ uc = 9.553344800e-11 luc = -1.889580518e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.182978791e-02 lu0 = -2.460846126e-09 wu0 = 3.388131789e-21
+ a0 = 1.962163306e+00 la0 = -1.889822803e-7
+ keta = -3.300858090e-01 lketa = 1.571043408e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.894409841e+00 lags = -1.828794488e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.165654879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 9.883424696e-10
+ nfactor = {1.180690296e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 5.151409622e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.224485132e-04 leta0 = -4.390393260e-10
+ etab = -8.696720778e-04 letab = 3.838919603e-10
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.674625680e-01 lpclm = 1.033798773e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.406254296e-02 lpdiblc2 = -1.986588152e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.847173507e-06 lalpha0 = 5.558777898e-11
+ alpha1 = 0.0
+ beta0 = 1.866091807e+01 lbeta0 = 2.512491472e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.633348340e-01 lkt1 = -1.059067758e-9
+ kt2 = -3.677703950e-02 lkt2 = 1.119453200e-9
+ at = 9.611513100e+04 lat = -2.182236985e-2
+ ute = -1.294833580e+00 lute = 1.190986724e-7
+ ua1 = 1.959366800e-09 lua1 = 2.118135515e-16
+ ub1 = -1.783685070e-18 lub1 = -3.666789859e-25
+ uc1 = -3.004568360e-11 luc1 = 1.898889909e-18 wuc1 = 3.155443621e-30
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.21 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {8.283814936e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.636354417e-07 wvth0 = 2.045122722e-06 pvth0 = -9.733761593e-13
+ k1 = 3.018764880e-01 lk1 = 6.763892604e-8
+ k2 = 3.299633297e-02 lk2 = -3.158792907e-08 wk2 = -1.158232344e-07 pk2 = 5.512606839e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.100012282e+04 lvsat = 5.077343083e-02 wvsat = 6.611892934e-01 pvsat = -3.146930442e-7
+ ua = -1.260293671e-09 lua = -1.707529780e-16 wua = -1.456011152e-15 pua = 6.929885079e-22
+ ub = 3.030780406e-18 lub = -2.132305529e-25 wub = -1.828317362e-24 pub = 8.701876484e-31
+ uc = 5.022947588e-11 luc = 2.666620352e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.911308685e-02 lu0 = -1.167832258e-09 wu0 = -3.844383695e-09 pu0 = 1.829734420e-15
+ a0 = 1.672471440e+00 la0 = -5.110343687e-8
+ keta = 3.197985042e-02 lketa = -1.522080981e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.899950380e-02 lags = -2.236893788e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.168740301e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.135193164e-9
+ nfactor = {-8.900210773e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 5.313145826e-06 wnfactor = 5.417898882e-05 pnfactor = -2.578648973e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -3.240309672e-03 leta0 = 1.542225543e-9
+ etab = 5.071496219e-02 letab = -2.416781472e-08 wetab = 5.691002614e-22 petab = 5.790239044e-28
+ dsub = 1.596959656e+00 ldsub = -2.841229483e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.776113220e-01 lpclm = 3.359577794e-9
+ pdiblc1 = 0.39
+ pdiblc2 = 5.344835880e-03 lpdiblc2 = 2.162604533e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.438650175e-03 lalpha0 = 7.416684422e-10 walpha0 = -1.323488980e-23 palpha0 = 1.262177448e-29
+ alpha1 = 0.0
+ beta0 = 1.801339785e+01 lbeta0 = 2.820678717e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.835456200e-01 lkt1 = 8.560255839e-9
+ kt2 = -4.209283920e-02 lkt2 = 3.649508067e-9
+ at = 5.171740660e+04 lat = -6.912729213e-4
+ ute = -1.230023608e+00 lute = 8.825236623e-8
+ ua1 = 2.284556120e-09 lua1 = 5.703969469e-17
+ ub1 = -2.723020220e-18 lub1 = 8.039757871e-26
+ uc1 = -4.960541280e-11 luc1 = 1.120834302e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.22 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {2.068711234e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -2.850725818e-07 wvth0 = -7.304009720e-06 pvth0 = 1.139060316e-12
+ k1 = 3.731197071e-01 lk1 = 5.154152067e-8
+ k2 = -1.039225143e-01 lk2 = -6.511155385e-10 wk2 = 4.136544084e-07 pk2 = -6.450940499e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.097935655e+05 lvsat = -6.870744754e-02 wvsat = -2.361390334e+00 pvsat = 3.682588225e-7
+ ua = -1.102040912e-09 lua = -2.065101890e-16 wua = 5.200039829e-15 pua = -8.109462114e-22
+ ub = 4.569362703e-19 lub = 3.683295296e-25 wub = 6.529704864e-24 pub = -1.018307474e-30
+ uc = 1.206245854e-10 luc = -1.323915464e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.374229402e-02 lu0 = -4.473301617e-09 wu0 = 1.372994177e-08 pu0 = -2.141184419e-15
+ a0 = 4.668449786e+00 la0 = -7.280447441e-7
+ keta = 7.382337983e-02 lketa = -2.467535528e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.655382929e+00 lags = 5.999837727e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.598193535e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.083868898e-8
+ nfactor = {4.035456925e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -5.815971721e-06 wnfactor = -1.934963886e-04 pnfactor = 3.017576181e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 7.038215705e-06 lcit = -4.605348385e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.910912508e-01 leta0 = 4.398714563e-08 weta0 = -2.541098842e-21 peta0 = 4.038967835e-28
+ etab = -1.436999391e-01 letab = 1.976023224e-8
+ dsub = 3.874366711e-01 ldsub = -1.083122984e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 9.611628143e-01 lpclm = -1.284938819e-7
+ pdiblc1 = -9.689896045e-01 lpdiblc1 = 3.070637011e-7
+ pdiblc2 = 2.556292929e-02 lpdiblc2 = -2.405673672e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.665019257e-03 lalpha0 = -1.855556660e-10
+ alpha1 = 0.0
+ beta0 = 3.073591653e+01 lbeta0 = -5.397437710e-8
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.046366429e-01 lkt1 = -3.186422755e-8
+ kt2 = -1.422247143e-02 lkt2 = -2.647801531e-9
+ at = -2.793795643e+04 lat = 1.730685636e-2
+ ute = 8.302498143e-01 lute = -3.772664135e-7
+ ua1 = 7.547183371e-09 lua1 = -1.132050933e-15
+ ub1 = -7.263227971e-18 lub1 = 1.106257520e-24
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.23 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 5.05e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-7.200396601e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 1.498331201e-07 wvth0 = 4.819566711e-06 pvth0 = -7.516114285e-13
+ k1 = 7.856554333e-01 lk1 = -1.279342583e-8
+ k2 = -2.870166058e-01 lk2 = 2.790240804e-08 wk2 = 6.775633855e-07 pk2 = -1.056660100e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.432375730e+05 lvsat = 4.051959494e-03 wvsat = 2.518799836e-01 pvsat = -3.928068345e-8
+ ua = -2.481319309e-09 lua = 8.588277042e-18 wua = 1.490992454e-15 pua = -2.325202732e-22
+ ub = -1.008738367e-17 lub = 2.012716225e-24 wub = 6.146453022e-23 pub = -9.585393487e-30
+ uc = 9.910064333e-11 luc = -9.882495878e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -7.160220510e-03 lu0 = 3.464945524e-09 wu0 = 9.531155192e-08 pu0 = -1.486383652e-14
+ a0 = 0.0
+ keta = -1.440907387e-02 lketa = -1.091550412e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.404198333e-01 lags = 3.921833199e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.424396780e-03+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.370705452e-8
+ nfactor = {-5.006538961e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.285020864e-06 wnfactor = 2.603936517e-04 pnfactor = -4.060838998e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.441633553e-07 lcit = 5.989976254e-13
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.154381393e-01 leta0 = -1.941111276e-8
+ etab = -3.860582515e-02 letab = 3.370805159e-9
+ dsub = 5.614173009e-01 ldsub = -3.796350905e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -4.137692667e-01 lpclm = 8.592677614e-8
+ pdiblc1 = 1.472992513e+00 lpdiblc1 = -7.376341016e-8
+ pdiblc2 = 4.039438833e-02 lpdiblc2 = -4.718639711e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.953879925e-03 lalpha0 = -5.425034872e-10
+ alpha1 = 0.0
+ beta0 = 3.551452838e+01 lbeta0 = -7.991988951e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.460355833e-01 lkt1 = 2.137693722e-8
+ kt2 = -1.120399083e-01 lkt2 = 1.260682775e-8
+ at = 1.189851300e+05 lat = -5.605798973e-3
+ ute = -2.280785333e+00 lute = 1.078995177e-7
+ ua1 = -6.950037167e-10 lua1 = 1.533181436e-16
+ ub1 = 1.068612467e-18 lub1 = -1.930929962e-25
+ uc1 = 1.083841733e-10 luc1 = -1.690251183e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.24 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.283833188e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 7.148930074e-10
+ k1 = 2.460777990e-01 wk1 = 7.631409306e-7
+ k2 = 5.176336310e-02 wk2 = -2.983889129e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.516973769e+05 wvsat = -5.380820208e-1
+ ua = -1.510533829e-09 wua = 1.211372227e-15
+ ub = 2.943208332e-18 wub = -1.396762665e-24
+ uc = 7.256765782e-11 wuc = -1.052270287e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.202014166e-02 wu0 = 1.871077995e-9
+ a0 = 2.282443201e+00 wa0 = -1.769730879e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.657893055e-01 wags = -9.036188775e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.249964441e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = 3.014833258e-8
+ nfactor = {5.563037292e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 2.301913561e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.743216080e-05 wcit = -3.677433166e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.271000965e-01 wpclm = 9.675620854e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.401939196e-03 wpdiblc2 = 9.156808583e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.630730053e-05 walpha0 = 3.702413969e-11
+ alpha1 = 0.0
+ beta0 = 1.716321658e+01 wbeta0 = 1.871033866e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.513990151e-01 wkt1 = -1.301811341e-8
+ kt2 = -3.455622111e-02 wkt2 = -6.619379698e-10
+ at = -3.040853166e+05 wat = 1.841548206e+0
+ ute = -1.101619698e+00 wute = -4.714469319e-7
+ ua1 = 4.174497588e-09 wua1 = -6.181029665e-15
+ ub1 = -5.033630251e-18 wub1 = 8.711103683e-24
+ uc1 = 2.518759799e-12 wuc1 = -1.459499675e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.25 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.283833188e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 7.148930074e-10
+ k1 = 2.460777990e-01 wk1 = 7.631409306e-7
+ k2 = 5.176336310e-02 wk2 = -2.983889129e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.516973769e+05 wvsat = -5.380820208e-1
+ ua = -1.510533829e-09 wua = 1.211372227e-15
+ ub = 2.943208332e-18 wub = -1.396762665e-24
+ uc = 7.256765782e-11 wuc = -1.052270287e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.202014166e-02 wu0 = 1.871077995e-9
+ a0 = 2.282443201e+00 wa0 = -1.769730879e-6
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.657893055e-01 wags = -9.036188775e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.249964441e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = 3.014833258e-8
+ nfactor = {5.563037292e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 2.301913561e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.743216080e-05 wcit = -3.677433166e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.271000965e-01 wpclm = 9.675620854e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 6.401939196e-03 wpdiblc2 = 9.156808583e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.630730053e-05 walpha0 = 3.702413969e-11
+ alpha1 = 0.0
+ beta0 = 1.716321658e+01 wbeta0 = 1.871033866e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.513990151e-01 wkt1 = -1.301811341e-8
+ kt2 = -3.455622111e-02 wkt2 = -6.619379698e-10
+ at = -3.040853166e+05 wat = 1.841548206e+0
+ ute = -1.101619698e+00 wute = -4.714469319e-7
+ ua1 = 4.174497588e-09 wua1 = -6.181029665e-15
+ ub1 = -5.033630251e-18 wub1 = 8.711103683e-24
+ uc1 = 2.518759799e-12 wuc1 = -1.459499675e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.26 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.427468825e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -5.710881119e-08 wvth0 = -6.164446835e-08 pvth0 = 2.479377028e-13
+ k1 = -7.769216345e-02 lk1 = 1.287293182e-06 wk1 = 1.900844946e-06 pk1 = -4.523454281e-12
+ k2 = 1.760949443e-01 lk2 = -4.943361503e-07 wk2 = -7.490101701e-07 pk2 = 1.791647588e-12
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.357099375e+05 lvsat = -1.129219740e+00 wvsat = -9.933743534e-01 pvsat = 1.810219550e-6
+ ua = -1.742434036e-09 lua = 9.220236246e-16 wua = 2.290298938e-15 pua = -4.289758656e-21
+ ub = 3.181789241e-18 lub = -9.485857673e-25 wub = -2.494792005e-24 pub = 4.365709756e-30
+ uc = 3.822578635e-11 luc = 1.365415639e-16 wuc = 3.289626637e-17 puc = -1.726316508e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.031056843e-02 lu0 = 6.797177696e-09 wu0 = 8.163365249e-09 pu0 = -2.501781951e-14
+ a0 = 2.526383963e+00 la0 = -9.698962734e-07 wa0 = -2.955223259e-06 pa0 = 4.713458429e-12
+ keta = 1.608135447e-01 lketa = -6.393866130e-07 wketa = 2.602106457e-07 pketa = -1.034584517e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.925508546e-01 lags = 1.086382419e-06 wags = -2.906420935e-06 pags = 1.119650997e-11
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.481005449e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 9.186074979e-08 wvoff = 1.075455585e-07 pvoff = -3.077275005e-13
+ nfactor = {-7.531616644e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 5.206368932e-06 wnfactor = 6.234323511e-06 pnfactor = -1.563506534e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.971482487e-05 lcit = -4.883525821e-11 wcit = -7.310645198e-11 pcit = 1.444546938e-16
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386527637e-01 letab = 2.729599558e-07 wetab = -5.689610042e-11 petab = 2.262160505e-16
+ dsub = 5.837108483e-01 ldsub = -9.427314735e-08 wdsub = 5.604374161e-07 pdsub = -2.228271145e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.039314373e-01 lpclm = -9.211743039e-08 wpclm = 9.464894556e-07 ppclm = 8.378372240e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 2.873828640e-03 lpdiblc2 = 1.402759117e-08 wpdiblc2 = 7.635669833e-09 ppdiblc2 = -2.671834016e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -5.628350342e-05 lalpha0 = 3.283769070e-10 walpha0 = -2.023117640e-11 palpha0 = 2.276442740e-16
+ alpha1 = 0.0
+ beta0 = 1.328208851e+01 lbeta0 = 1.543117114e-05 wbeta0 = 2.615638872e-06 pbeta0 = -2.960512276e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.219970379e-01 lkt1 = -1.169007910e-07 wkt1 = -1.068276481e-07 pkt1 = 3.729820194e-13
+ kt2 = -6.825592126e-02 lkt2 = 1.339883228e-07 wkt2 = 1.033060575e-07 pkt2 = -4.133715517e-13
+ at = -6.848108433e+05 lat = 1.513745658e+00 wat = 3.773603168e+00 pat = -7.681753924e-6
+ ute = -9.375003696e-01 lute = -6.525302457e-07 wute = -1.105079110e-06 pute = 2.519289860e-12
+ ua1 = 5.111926099e-09 lua1 = -3.727168888e-15 wua1 = -9.373896399e-15 pua1 = 1.269467849e-20
+ ub1 = -6.613924960e-18 lub1 = 6.283172746e-24 wub1 = 1.458673418e-23 pub1 = -2.336121308e-29
+ uc1 = 2.349053789e-11 luc1 = -8.338274110e-17 wuc1 = -1.885094132e-16 puc1 = 1.692142283e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.27 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.986365752e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 3.005095053e-08 wvth0 = 1.036120486e-07 pvth0 = -7.860091188e-14
+ k1 = 7.117532471e-01 lk1 = -2.726114768e-07 wk1 = -7.827688109e-07 pk1 = 7.792323222e-13
+ k2 = -1.222754883e-01 lk2 = 9.522890597e-08 wk2 = 3.116351996e-07 pk2 = -3.041346307e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.072640805e+04 lvsat = 6.918964658e-03 wvsat = -1.824630183e-01 pvsat = 2.078992970e-7
+ ua = -9.627034924e-10 lua = -6.186849421e-16 wua = -7.641820989e-17 pua = 3.867560920e-22
+ ub = 2.536055133e-18 lub = 3.273525432e-25 wub = 8.975251501e-26 pub = -7.412209894e-31
+ uc = 1.338908825e-10 luc = -5.248788286e-17 wuc = -8.861579946e-17 puc = 6.747011570e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.673113121e-02 lu0 = -5.889533334e-09 wu0 = -2.183972524e-09 pu0 = -4.571997435e-15
+ a0 = 1.981708690e+00 la0 = 1.063548320e-07 wa0 = 4.297977374e-07 pa0 = -1.975173808e-12
+ keta = -1.802883527e-01 lketa = 3.461368119e-08 wketa = -4.031330689e-07 pketa = 2.761494961e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.346473899e-01 lags = 2.128099790e-06 wags = 5.093060565e-06 pags = -4.610065501e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.879879364e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.531654566e-08 wvoff = -9.129405759e-08 pvoff = 8.516963895e-14
+ nfactor = {2.260684036e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -7.488394797e-07 wnfactor = -4.355238607e-06 pnfactor = 5.289379929e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.169151556e-04 leta0 = -3.342350169e-11 weta0 = 4.866671658e-11 peta0 = -9.616299863e-17
+ etab = -5.409291714e-04 letab = 5.787638084e-11 wetab = 8.816680583e-11 petab = -6.042099914e-17
+ dsub = -2.283463502e-01 ldsub = 1.510311274e-06 wdsub = 4.204600898e-07 pdsub = -1.951682947e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.302785382e-01 lpclm = 1.343108124e-06 wpclm = 3.270082525e-06 ppclm = -4.507520002e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.710653061e-03 lpdiblc2 = 5.183679504e-10 wpdiblc2 = -2.025139449e-08 ppdiblc2 = 2.838510459e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.406117439e-04 lalpha0 = -6.067825705e-11 walpha0 = 2.776493280e-10 palpha0 = -3.609527086e-16
+ alpha1 = 0.0
+ beta0 = 2.033771694e+01 lbeta0 = 1.489602139e-06 wbeta0 = 5.243865712e-06 pbeta0 = -8.153757100e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.986121654e-01 lkt1 = 3.448687006e-08 wkt1 = 1.674229741e-07 pkt1 = -1.689234976e-13
+ kt2 = 5.519006838e-02 lkt2 = -1.099347804e-07 wkt2 = -3.146310761e-07 pkt2 = 4.124513274e-13
+ at = 9.351288859e+04 lat = -2.418312012e-02 wat = -2.495499670e-01 pat = 2.677955128e-7
+ ute = -1.263919490e+00 lute = -7.542383891e-09 wute = -1.416269977e-07 pute = 6.155566579e-13
+ ua1 = 5.008681497e-09 lua1 = -3.523162717e-15 wua1 = -9.583192175e-15 pua1 = 1.310823648e-20
+ ub1 = -5.984196174e-18 lub1 = 5.038860151e-24 wub1 = 1.192378134e-23 pub1 = -1.809935141e-29
+ uc1 = -9.618303716e-11 luc1 = 1.530862595e-16 wuc1 = 2.254268380e-16 puc1 = -6.487031074e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.28 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.355386013e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -5.963581852e-09 wvth0 = 2.790614879e-08 pvth0 = -4.715738964e-15
+ k1 = 4.029067816e-01 lk1 = 2.880723122e-08 wk1 = 1.221525546e-07 pk1 = -1.039256845e-13
+ k2 = -7.877157950e-03 lk2 = -1.641814451e-08 wk2 = -4.238251851e-08 pk2 = 4.136896133e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -7.261414148e+04 lvsat = 1.370526740e-01 wvsat = 1.899450496e-01 pvsat = -1.555523568e-7
+ ua = -1.063872918e-09 lua = -5.199486407e-16 wua = -1.906146817e-15 pua = 2.172479726e-21
+ ub = 2.600905729e-18 lub = 2.640616038e-25 wub = 1.391318895e-24 pub = -2.011484698e-30
+ uc = 9.264506714e-11 luc = -1.223402937e-17 wuc = 1.429170850e-17 puc = -3.296246669e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.701065640e-02 lu0 = -6.162335949e-09 wu0 = -2.563493730e-08 pu0 = 1.831497164e-14
+ a0 = 2.932411928e+00 la0 = -8.214839925e-07 wa0 = -4.800790182e-06 pa0 = 3.129618472e-12
+ keta = -2.998023213e-01 lketa = 1.512533388e-07 wketa = -1.498426970e-07 pketa = 2.895075762e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.818607252e+00 lags = -2.803624077e-06 wags = -4.572928788e-06 pags = 4.823456809e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.102363468e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -4.394565621e-09 wvoff = -3.131658977e-08 pvoff = 2.663462923e-14
+ nfactor = {1.075685707e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 4.076596392e-07 wnfactor = 5.195627065e-07 pnfactor = 5.318175864e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 9.562691322e-04 leta0 = -4.622109218e-10 weta0 = -1.673444058e-10 peta0 = 1.146530562e-16
+ etab = -9.313929843e-04 letab = 4.389495390e-10 wetab = 3.053950453e-10 petab = -2.724248994e-16
+ dsub = 1.623013307e+00 ldsub = -2.965231836e-07 wdsub = -3.082669844e-06 pdsub = 1.467196712e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.713482997e-01 lpclm = -2.480958890e-08 wpclm = -1.998426601e-06 ppclm = 6.342814785e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.203170526e-02 lpdiblc2 = -1.746862941e-09 wpdiblc2 = 1.004858495e-08 ppdiblc2 = -1.186160343e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.507539435e-05 lalpha0 = 5.207944333e-11 walpha0 = -1.099852367e-10 palpha0 = 1.735924481e-17
+ alpha1 = 0.0
+ beta0 = 1.961327591e+01 lbeta0 = 2.196620365e-06 wbeta0 = -4.712266608e-06 pbeta0 = 1.562930238e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.509415498e-01 lkt1 = -1.203726722e-08 wkt1 = -6.132197030e-08 pkt1 = 5.432013093e-14
+ kt2 = -6.592878368e-02 lkt2 = 8.271163264e-09 wkt2 = 1.442428302e-07 pkt2 = -3.538666140e-14
+ at = 1.168712449e+05 lat = -4.697970793e-02 wat = -1.027012514e-01 pat = 1.244785088e-7
+ ute = -2.191987518e+00 lute = 8.982056077e-07 wute = 4.439117686e-06 pute = -3.855021116e-12
+ ua1 = -2.543334240e-09 lua1 = 3.847227042e-15 wua1 = 2.227936475e-14 pua1 = -1.798802595e-20
+ ub1 = 4.348914792e-18 lub1 = -5.045739496e-24 wub1 = -3.034410412e-23 pub1 = 2.315199140e-29
+ uc1 = 1.801030957e-10 luc1 = -1.165551918e-16 wuc1 = -1.039816160e-15 puc1 = 5.861107964e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.29 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.968637400e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.515128160e-08 wvth0 = -3.475900900e-09 pvth0 = 1.022054759e-14
+ k1 = 3.240912574e-01 lk1 = 6.631947994e-08 wk1 = -1.099186792e-07 pk1 = 6.528619293e-15
+ k2 = -7.976668176e-04 lk2 = -1.978762831e-08 wk2 = 5.138947659e-08 pk2 = -3.261819739e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.733382112e+05 lvsat = -2.760334829e-02 wvsat = -2.904995679e-01 pvsat = 7.311525887e-8
+ ua = -3.095069079e-09 lua = 4.467991719e-16 wua = 7.622457566e-15 pua = -2.362659530e-21
+ ub = 4.078275261e-18 lub = -4.390924245e-25 wub = -7.011321901e-24 pub = 1.987752189e-30
+ uc = 5.186234121e-11 luc = 7.176509034e-18 wuc = -8.079417652e-18 puc = -2.231492920e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.727173645e-02 lu0 = 3.232403002e-09 wu0 = 5.474661809e-08 pu0 = -1.994262965e-14
+ a0 = 1.054428248e+00 la0 = 7.234234001e-08 wa0 = 3.058077715e-06 pa0 = -6.108097040e-13
+ keta = 6.911682585e-02 lketa = -2.433372925e-08 wketa = -1.837537544e-07 pketa = 4.509072538e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.040831824e+00 lags = 4.611259505e-07 wags = 1.058788541e-05 pags = -2.392332708e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.248181020e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.545620772e-09 wvoff = 3.930726785e-08 pvoff = -6.978795805e-15
+ nfactor = {1.402066072e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.523189045e-07 wnfactor = 3.203322989e-06 pnfactor = -7.455181202e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.940011850e-03 leta0 = -1.406373174e-09 weta0 = -3.058023104e-08 peta0 = 1.458966645e-14
+ etab = 1.013801562e-01 letab = -4.825623229e-08 wetab = -2.506913799e-07 petab = 1.191894902e-13
+ dsub = 1.495761755e+00 ldsub = -2.359578074e-07 wdsub = 5.007272125e-07 pdsub = -2.383211168e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 5.932494683e-01 lpclm = -3.523345009e-08 wpclm = -1.066977548e-06 ppclm = 1.909583019e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 5.367464848e-03 lpdiblc2 = 1.424982282e-09 wpdiblc2 = -1.119681315e-10 ppdiblc2 = 3.649754895e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.187419176e-03 lalpha0 = 6.291662339e-10 walpha0 = -1.243090987e-09 palpha0 = 5.566609267e-16
+ alpha1 = 0.0
+ beta0 = 1.852664409e+01 lbeta0 = 2.713802778e-06 wbeta0 = -2.539542396e-06 pbeta0 = 5.288221491e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.379202211e-01 lkt1 = 2.936023140e-08 wkt1 = 2.690455263e-07 pkt1 = -1.029182791e-13
+ kt2 = -5.908798628e-02 lkt2 = 5.015285743e-09 wkt2 = 8.409198776e-08 pkt2 = -6.757867940e-15
+ at = 9.910017228e+02 lat = 8.173493792e-03 wat = 2.509942513e-01 pat = -4.386286570e-8
+ ute = -9.665554815e-01 lute = 3.149612299e-07 wute = -1.303640290e-06 pute = -1.121755457e-12
+ ua1 = 4.863232633e-09 lua1 = 3.220715382e-16 wua1 = -1.275929139e-14 pua1 = -1.311377562e-21
+ ub1 = -6.499755974e-18 lub1 = 1.176853554e-25 wub1 = 1.868728851e-23 pub1 = -1.844999189e-31
+ uc1 = -1.638464744e-10 luc1 = 4.714760605e-17 wuc1 = 5.652647727e-16 puc1 = -1.778274735e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.30 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.288088727e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -6.496428433e-08 wvth0 = -1.793728345e-07 pvth0 = 4.996445974e-14
+ k1 = 3.888208930e-01 lk1 = 5.169381879e-08 wk1 = -7.768946746e-08 pk1 = -7.535711079e-16
+ k2 = -2.979173862e-02 lk2 = -1.323641779e-08 wk2 = 4.685533055e-08 pk2 = -2.237329443e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.308715321e+04 lvsat = 1.312437827e-02 wvsat = 1.952729942e-01 pvsat = -3.664505154e-8
+ ua = 2.394361061e-09 lua = -7.935375682e-16 wua = -1.210015713e-14 pua = 2.093665261e-21
+ ub = 6.340580361e-20 lub = 4.680673293e-25 wub = 8.476893613e-24 pub = -1.511810106e-30
+ uc = 2.011244503e-10 luc = -2.654926451e-17 wuc = -3.983133314e-16 puc = 6.585842361e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 7.261993500e-02 lu0 = -9.273522459e-09 wu0 = -1.291566258e-07 pu0 = 2.161030831e-14
+ a0 = 4.437005751e+00 la0 = -6.919510469e-07 wa0 = 1.145185082e-06 pa0 = -1.785916136e-13
+ keta = -2.450350375e-02 lketa = -3.180215773e-09 wketa = 4.865214200e-07 pketa = -1.063579503e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.822285477e+00 lags = 6.376954036e-07 wags = 8.258338112e-07 pags = -1.865971496e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.722597243e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.326505532e-08 wvoff = 6.155495452e-08 pvoff = -1.200566061e-14
+ nfactor = {1.127102009e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.144470347e-07 wnfactor = 6.011192857e-07 pnfactor = -1.575501933e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.006788508e-05 lcit = -1.145088634e-12 wcit = -1.499080406e-11 pcit = 3.387172178e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.489989820e-01 leta0 = 5.551924241e-08 weta0 = 2.865274535e-07 peta0 = -5.706081488e-14
+ etab = -3.170663457e-01 letab = 4.629175481e-08 wetab = 8.578169796e-07 petab = -1.312779737e-13
+ dsub = 8.066516601e-01 ldsub = -8.025338143e-08 wdsub = -2.074275765e-06 pdsub = 3.435008061e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.351136998e+00 lpclm = -2.064781375e-07 wpclm = -1.929592263e-06 ppclm = 3.858660969e-13
+ pdiblc1 = -9.788240722e-01 lpdiblc1 = 3.092857991e-07 wpdiblc1 = 4.866094648e-08 ppdiblc1 = -1.099494086e-14
+ pdiblc2 = 2.230777451e-02 lpdiblc2 = -2.402680686e-09 wpdiblc2 = 1.610650584e-08 ppdiblc2 = -1.480929759e-17
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.212332501e-03 lalpha0 = 6.347953998e-10 walpha0 = 1.918513650e-08 palpha0 = -4.059097074e-15
+ alpha1 = 0.0
+ beta0 = 2.510144258e+01 lbeta0 = 1.228227059e-06 wbeta0 = 2.787937708e-05 pbeta0 = -6.344332706e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 3.848443528e-02 lkt1 = -5.568840071e-08 wkt1 = -7.081630946e-07 pkt1 = 1.178820088e-13
+ kt2 = -1.855983482e-02 lkt2 = -4.142050080e-09 wkt2 = 2.146127406e-08 pkt2 = 7.393541822e-15
+ at = -1.067450997e+05 lat = 3.251646590e-02 wat = 3.899377447e-01 pat = -7.525714803e-8
+ ute = 4.472987254e+00 lute = -9.141034512e-07 wute = -1.802426485e-05 pute = 2.656269662e-12
+ ua1 = 1.862035468e-08 lua1 = -2.786350188e-15 wua1 = -5.479005162e-14 pua1 = 8.185472713e-21
+ ub1 = -1.759539402e-17 lub1 = 2.624744771e-24 wub1 = 5.112355759e-23 pub1 = -7.513474918e-30
+ uc1 = 1.248690445e-10 luc1 = -1.808766544e-17 wuc1 = -6.178520321e-16 puc1 = 8.949776859e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.31 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.01e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.119889890e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 1.563377653e-08 wvth0 = 7.026889552e-07 pvth0 = -8.759307636e-14
+ k1 = 6.486287589e-01 lk1 = 1.117678210e-08 wk1 = 6.780079850e-07 pk1 = -1.186045888e-13
+ k2 = -1.035597703e-01 lk2 = -1.732293258e-09 wk2 = -2.301810370e-07 pk2 = 4.096649208e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.375108407e+05 lvsat = -9.398495797e-03 wvsat = -2.145841450e-01 pvsat = 2.727216933e-8
+ ua = -2.926540194e-09 lua = 3.625698244e-17 wua = 3.693945393e-15 pua = -3.694250275e-22
+ ub = 1.539373030e-18 lub = 2.378902404e-25 wub = 3.935338051e-24 pub = -8.035545163e-31
+ uc = 1.186074377e-10 luc = -1.368073639e-17 wuc = -9.651961831e-17 puc = 1.879369406e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.094064550e-02 lu0 = 3.757750069e-09 wu0 = 1.140170948e-07 pu0 = -1.631263341e-14
+ a0 = 0.0
+ keta = -2.760936010e-01 lketa = 3.605525989e-08 wketa = 1.294815040e-06 pketa = -2.324113403e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.302400748e+00 lags = -5.549413224e-09 wags = -1.791081565e-06 pags = 2.215108033e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {1.940799623e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -4.386561881e-08 wvoff = -9.723035690e-07 pvoff = 1.492245761e-13
+ nfactor = {5.180685673e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -3.177093378e-07 wnfactor = -1.296392885e-05 pnfactor = 1.957919063e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.437762326e-05 lcit = -3.376692303e-12 wcit = -1.194123596e-10 pcit = 1.967171376e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.100160203e-01 leta0 = -4.725414719e-08 weta0 = -9.627713551e-07 peta0 = 1.377673343e-13
+ etab = 1.846722419e-02 letab = -6.034705415e-09 wetab = -2.823974481e-07 petab = 4.653846632e-14
+ dsub = 4.265648323e-01 ldsub = -2.097884062e-08 wdsub = 6.672500149e-07 pdsub = -8.404013938e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.612890665e+00 lpclm = 2.557619765e-07 wpclm = 5.933252677e-06 ppclm = -8.403445715e-13
+ pdiblc1 = 2.199022170e+00 lpdiblc1 = -1.862993224e-07 wpdiblc1 = -3.592394741e-06 ppdiblc1 = 5.568276936e-13
+ pdiblc2 = 4.169342426e-02 lpdiblc2 = -5.425872764e-09 wpdiblc2 = -6.427629753e-09 ppdiblc2 = 3.499389147e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.019452451e-02 lalpha0 = -1.144103951e-09 walpha0 = -2.593070940e-08 palpha0 = 2.976719094e-15
+ alpha1 = 0.0
+ beta0 = 4.143977481e+01 lbeta0 = -1.319735853e-06 wbeta0 = -2.931811938e-05 pbeta0 = 2.575616866e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -9.919943370e-01 lkt1 = 1.050147638e-07 wkt1 = 2.701403913e-06 pkt1 = -4.138399660e-13
+ kt2 = -1.825480548e-01 lkt2 = 2.143191283e-08 wkt2 = 3.488743089e-07 pkt2 = -4.366652097e-14
+ at = 2.949994955e+05 lat = -3.013560372e-02 wat = -8.709190805e-01 pat = 1.213734739e-7
+ ute = -2.732550466e+00 lute = 2.096001563e-07 wute = 2.235333879e-06 pute = -5.032147597e-13
+ ua1 = -5.809072749e-10 lua1 = 2.080866138e-16 wua1 = -5.645491938e-16 pua1 = -2.709943906e-22
+ ub1 = 3.773868161e-19 lub1 = -1.781103997e-25 wub1 = 3.420184519e-24 pub1 = -7.413388733e-32
+ uc1 = 7.099962758e-11 luc1 = -9.686729872e-18 wuc1 = 1.849787324e-16 puc1 = -3.570368913e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.32 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.428625+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.50407
+ k2 = -0.049111861
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.10100975e-9
+ ub = 2.47101e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03265269
+ a0 = 1.6841569
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.535241
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11480431+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.33450304+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.33 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.428625+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.50407
+ k2 = -0.049111861
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 169790.0
+ ua = -1.10100975e-9
+ ub = 2.47101e-18
+ uc = 6.9010287e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.03265269
+ a0 = 1.6841569
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.535241
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11480431+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.33450304+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.2558
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.34 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.219069676e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 2.671056094e-8
+ k1 = 5.649193802e-01 lk1 = -2.419340934e-7
+ k2 = -7.712012334e-02 lk2 = 1.113594506e-07 wk2 = -1.355252716e-20
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.998835841e+05 lvsat = -5.172455856e-1
+ ua = -9.681612372e-10 lua = -5.281990446e-16
+ ub = 2.338384236e-18 lub = 5.273134064e-25
+ uc = 4.934690412e-11 luc = 7.818062715e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.307032679e-02 lu0 = -1.660503003e-9
+ a0 = 1.527322686e+00 la0 = 6.235649940e-7
+ keta = 2.487819847e-01 lketa = -9.891447323e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.900120038e-01 lags = 4.871544681e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.117430201e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.217153572e-8
+ nfactor = {1.354452775e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -7.931914723e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386719983e-01 letab = 2.730364318e-7
+ dsub = 7.731758301e-01 ldsub = -8.475764417e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.160447140e-01 lpclm = -6.379298063e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 5.455190990e-03 lpdiblc2 = 4.995021808e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -6.312298158e-05 lalpha0 = 4.053357555e-10 palpha0 = 2.524354897e-29
+ alpha1 = 0.0
+ beta0 = 1.416634776e+01 lbeta0 = 1.443032182e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.581118615e-01 lkt1 = 9.191845731e-9
+ kt2 = -3.333162865e-02 lkt2 = -5.758652069e-9
+ at = 5.909170702e+05 lat = -1.083196169e+0
+ ute = -1.311090332e+00 lute = 1.991566575e-7
+ ua1 = 1.942927992e-09 lua1 = 5.644736032e-16
+ ub1 = -1.682642275e-18 lub1 = -1.614465212e-24
+ uc1 = -4.023813460e-11 luc1 = -2.617711964e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.35 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.336643131e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 3.478634142e-9
+ k1 = 4.471255220e-01 lk1 = -9.179319196e-9
+ k2 = -1.692214156e-02 lk2 = -7.588751450e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -9.581823000e+02 lvsat = 7.720270267e-2
+ ua = -9.885379109e-10 lua = -4.879357562e-16
+ ub = 2.566397431e-18 lub = 7.677073470e-26
+ uc = 1.039328705e-10 luc = -2.967851311e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.599280378e-02 lu0 = -7.435171412e-9
+ a0 = 2.127008804e+00 la0 = -5.613847923e-7
+ keta = -3.165740420e-01 lketa = 1.279705088e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.487144552e+00 lags = 5.695921835e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.196622343e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.476435734e-9
+ nfactor = {7.883248042e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.039321416e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.333677305e-04 leta0 = -6.593296708e-11
+ etab = -5.111229490e-04 letab = 3.745007958e-11
+ dsub = -8.620297978e-02 ldsub = 8.505131177e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.752260340e-01 lpclm = -1.807323099e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.864339845e-03 lpdiblc2 = 1.011441413e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.344756141e-04 lalpha0 = -1.827041896e-10
+ alpha1 = 0.0
+ beta0 = 2.211049102e+01 lbeta0 = -1.266908037e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.420121065e-01 lkt1 = -2.262046516e-8
+ kt2 = -5.117608310e-02 lkt2 = 2.950109770e-8
+ at = 9.148464300e+03 lat = 6.634950762e-2
+ ute = -1.311798800e+00 lute = 2.005565539e-7
+ ua1 = 1.768927550e-09 lua1 = 9.082897776e-16
+ ub1 = -1.953168000e-18 lub1 = -1.079919905e-24
+ uc1 = -1.997382890e-11 luc1 = -6.621837449e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.36 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.449727287e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -7.557814091e-9
+ k1 = 4.442024390e-01 lk1 = -6.326536342e-9
+ k2 = -2.220525752e-02 lk2 = -2.432694433e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -8.400128760e+03 lvsat = 8.446567031e-2
+ ua = -1.708276846e-09 lua = 2.144934575e-16
+ ub = 3.071263706e-18 lub = -4.159535069e-25
+ uc = 9.747661160e-11 luc = -2.337752724e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.834434900e-02 lu0 = 2.933803490e-11
+ a0 = 1.309426741e+00 la0 = 2.365344226e-7
+ keta = -3.504590816e-01 lketa = 1.610406132e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.272654315e+00 lags = -1.172976069e-06 wags = 4.336808690e-19 pags = -2.067951531e-25
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.208234292e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.609703896e-9
+ nfactor = {1.251332329e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 5.874492221e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.996955390e-04 leta0 = -4.234505918e-10
+ etab = -8.281492232e-04 letab = 3.468518719e-10
+ dsub = 5.808666392e-01 ldsub = 1.994865231e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.042523090e-01 lpclm = 1.896195790e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 1.542879280e-02 lpdiblc2 = -2.147863733e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.210690339e-05 lalpha0 = 5.794801832e-11
+ alpha1 = 0.0
+ beta0 = 1.802021756e+01 lbeta0 = 2.724994347e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.716724390e-01 lkt1 = 6.326536342e-9
+ kt2 = -1.716514940e-02 lkt2 = -3.691873043e-9
+ at = 8.215141680e+04 lat = -4.897723876e-3
+ ute = -6.912716000e-01 lute = -4.050469670e-7
+ ua1 = 4.988567297e-09 lua1 = -2.233917634e-15
+ ub1 = -5.909403030e-18 lub1 = 2.781167672e-24
+ uc1 = -1.714236656e-10 luc1 = 8.158909364e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.37 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.956886552e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.169605930e-8
+ k1 = 2.869314605e-01 lk1 = 6.852658585e-8
+ k2 = 1.657538139e-02 lk2 = -2.089033952e-08 pk2 = -1.615587134e-27
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.751301085e+05 lvsat = -2.885546099e-3
+ ua = -5.181733502e-10 lua = -3.519363013e-16
+ ub = 1.707983881e-18 lub = 2.328995259e-25
+ uc = 4.913096269e-11 luc = -3.674156442e-19
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.577972093e-02 lu0 = -3.509527236e-9
+ a0 = 2.088261147e+00 la0 = -1.341518128e-7
+ keta = 6.995881154e-03 lketa = -9.090076313e-09 pketa = 8.077935669e-28
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.538575008e+00 lags = -3.476410231e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.115296410e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.863253677e-10
+ nfactor = {2.485001498e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.843811626e-10
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -7.398132812e-03 leta0 = 3.525900812e-09 weta0 = -2.646977960e-23 peta0 = -1.104405267e-29
+ etab = 1.662985872e-02 letab = -7.962287009e-09 wetab = -4.499862532e-22 petab = 1.577721810e-28
+ dsub = 1.665040732e+00 ldsub = -3.165261363e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.325403581e-01 lpclm = 2.932310906e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 5.329612200e-03 lpdiblc2 = 2.658841273e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.607666298e-03 lalpha0 = 8.173545120e-10 walpha0 = 7.940933881e-23 palpha0 = -6.310887242e-30
+ alpha1 = 0.0
+ beta0 = 1.766811049e+01 lbeta0 = 2.892579704e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.469650060e-01 lkt1 = -5.432966394e-9
+ kt2 = -3.065932240e-02 lkt2 = 2.730678596e-9
+ at = 8.584368980e+04 lat = -6.655061210e-3
+ ute = -1.407272280e+00 lute = -6.426644333e-8
+ ua1 = 5.497467010e-10 lua1 = -1.212609708e-16
+ ub1 = -1.822142192e-19 lub1 = 5.531215763e-26
+ uc1 = 2.725047380e-11 luc1 = -1.296986301e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.38 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.681689692e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -4.807298624e-8
+ k1 = 3.625567052e-01 lk1 = 5.143906183e-8
+ k2 = -1.395153221e-02 lk2 = -1.399278339e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.591023643e+05 lvsat = 7.359227087e-4
+ ua = -1.696293818e-09 lua = -8.573998159e-17
+ ub = 2.929157532e-18 lub = -4.302466066e-26
+ uc = 6.646815162e-11 luc = -4.284753482e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.895643743e-02 lu0 = -1.967806330e-9
+ a0 = 4.824154190e+00 la0 = -7.523268460e-7
+ keta = 1.399729736e-01 lketa = -3.913625035e-08 pketa = 3.231174268e-27
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.543098929e+00 lags = 5.746132029e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.514500710e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 9.206346523e-9
+ nfactor = {1.330320158e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.611846299e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.521337171e-01 leta0 = 3.622890608e-08 weta0 = 1.016439537e-20 peta0 = 2.827277484e-27
+ etab = -2.706736678e-02 letab = 1.911101093e-9
+ dsub = 1.054090078e-01 ldsub = 3.587265173e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 6.988069568e-01 lpclm = -7.602982891e-8
+ pdiblc1 = -9.623734480e-01 lpdiblc1 = 3.055687806e-07 ppdiblc1 = -2.584939414e-26
+ pdiblc2 = 2.775284071e-02 lpdiblc2 = -2.407687209e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.273514862e-03 lalpha0 = -7.374483709e-10
+ alpha1 = 0.0
+ beta0 = 3.452651935e+01 lbeta0 = -9.165777774e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.009216143e-01 lkt1 = -1.583647075e-8
+ kt2 = -1.130450214e-02 lkt2 = -1.642543041e-9
+ at = 2.507969571e+04 lat = 7.074563253e-3
+ ute = -1.620408571e+00 lute = -1.610829829e-8
+ ua1 = 9.768678643e-11 lua1 = -1.911803314e-17 pua1 = 7.523163845e-37
+ ub1 = -3.122440529e-19 lub1 = 8.469239854e-26 pub1 = -5.605193857e-45
+ uc1 = -8.400588186e-11 luc1 = 1.216851056e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.39 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 3.01e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.430259409e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 4.195319193e-07 wvth0 = 8.222659715e-06 pvth0 = -1.282323783e-12
+ k1 = 8.778403833e-01 lk1 = -2.891942778e-8
+ k2 = 8.616071726e-01 lk2 = -1.505361634e-07 wk2 = -3.085144854e-06 pk2 = 4.811283400e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.473985752e+06 lvsat = -5.162201416e-01 wvsat = -9.788076932e+00 pvsat = 1.526450597e-6
+ ua = 2.881062127e-09 lua = -7.995786412e-16 wua = -1.348494227e-14 pua = 2.102976747e-21
+ ub = 1.525669878e-18 lub = 1.758492390e-25 wub = 3.975871973e-24 pub = -6.200372342e-31
+ uc = 8.597741118e-11 luc = -7.327222511e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -2.957560498e-02 lu0 = 7.160265685e-09 wu0 = 1.691393049e-07 pu0 = -2.637727460e-14
+ a0 = 0.0
+ keta = 1.616396783e-01 lketa = -4.251517295e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 6.968965000e-01 lags = 6.933591582e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.346230698e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 6.582175686e-9
+ nfactor = {-6.195178268e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.013002857e-05 wnfactor = 1.856139125e-04 pnfactor = -2.894648966e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.599166667e-05 lcit = 3.273650417e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 8.453550807e-02 leta0 = -6.796595860e-10
+ etab = -7.700182521e-02 letab = 9.698379886e-9
+ dsub = 6.521395499e-01 ldsub = -4.938997632e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.929418833e-01 lpclm = -2.833017071e-8
+ pdiblc1 = 9.845547120e-01 lpdiblc1 = 1.945334024e-9
+ pdiblc2 = 3.952045950e-02 lpdiblc2 = -4.242847359e-09 ppdiblc2 = 8.077935669e-28
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.428226537e-03 lalpha0 = -1.377756568e-10
+ alpha1 = 0.0
+ beta0 = 3.152830782e+01 lbeta0 = -4.490066891e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -7.874081667e-02 lkt1 = -3.489056614e-8
+ kt2 = -6.460542167e-02 lkt2 = 6.669735359e-9
+ at = 5.711383333e+02 lat = 1.089667278e-2
+ ute = -1.976859500e+00 lute = 3.948022403e-8
+ ua1 = -7.717623100e-10 lua1 = 1.164725534e-16 wua1 = -2.524354897e-29 pua1 = 6.018531076e-36
+ ub1 = 1.533635808e-18 lub1 = -2.031725658e-25
+ uc1 = 1.335346960e-10 luc1 = -2.175694256e-17 wuc1 = -3.155443621e-30 puc1 = 1.504632769e-36
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.40 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.353395593e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = -1.979452070e-8
+ k1 = 4.695176889e-01 wk1 = 1.018602132e-7
+ k2 = -3.928860344e-02 wk2 = -2.895896329e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.333792741e+05 wvsat = 1.073388200e-1
+ ua = -1.245108299e-09 wua = 4.248025229e-16
+ ub = 2.668593822e-18 wub = -5.824771079e-25
+ uc = 1.242415467e-10 wuc = -1.628217536e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.436466883e-02 wu0 = -5.046913590e-9
+ a0 = 1.404023239e+00 wa0 = 8.258340336e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.329505333e-01 wags = 6.752295733e-9
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.202140963e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = 1.594805013e-8
+ nfactor = {9.145169641e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 1.238118952e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -9.185185185e-07 wcit = 1.744779259e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.696355704e-03 wpdiblc2 = 2.992645385e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.537812311e-05 walpha0 = 1.015818860e-11
+ alpha1 = 0.0
+ beta0 = 1.779857550e+01 wbeta0 = -8.329576184e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.536338222e-01 wkt1 = -6.385892089e-9
+ kt2 = -3.290501333e-02 wkt2 = -5.527460693e-9
+ at = 6.265388889e+05 wat = -9.081576044e-1
+ ute = -1.355933037e+00 wute = 2.798625932e-7
+ ua1 = 2.228483259e-09 wua1 = -4.232834483e-16
+ ub1 = -2.825792296e-18 wub1 = 2.172948089e-24
+ uc1 = -1.773134963e-10 wuc1 = 3.846889311e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.41 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.353395593e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = -1.979452070e-8
+ k1 = 4.695176889e-01 wk1 = 1.018602132e-7
+ k2 = -3.928860344e-02 wk2 = -2.895896329e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.333792741e+05 wvsat = 1.073388200e-1
+ ua = -1.245108299e-09 wua = 4.248025229e-16
+ ub = 2.668593822e-18 wub = -5.824771079e-25
+ uc = 1.242415467e-10 wuc = -1.628217536e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.436466883e-02 wu0 = -5.046913590e-9
+ a0 = 1.404023239e+00 wa0 = 8.258340336e-7
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 5.329505333e-01 wags = 6.752295733e-9
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.202140963e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = 1.594805013e-8
+ nfactor = {9.145169641e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 1.238118952e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -9.185185185e-07 wcit = 1.744779259e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 5.696355704e-03 wpdiblc2 = 2.992645385e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.537812311e-05 walpha0 = 1.015818860e-11
+ alpha1 = 0.0
+ beta0 = 1.779857550e+01 wbeta0 = -8.329576184e-9
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.536338222e-01 wkt1 = -6.385892089e-9
+ kt2 = -3.290501333e-02 wkt2 = -5.527460693e-9
+ at = 6.265388889e+05 wat = -9.081576044e-1
+ ute = -1.355933037e+00 wute = 2.798625932e-7
+ ua1 = 2.228483259e-09 wua1 = -4.232834483e-16
+ ub1 = -2.825792296e-18 wub1 = 2.172948089e-24
+ uc1 = -1.773134963e-10 wuc1 = 3.846889311e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.42 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.335320130e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 7.186713400e-09 wvth0 = -3.427063396e-08 pvth0 = 5.755630255e-14
+ k1 = 5.142985559e-01 lk1 = -1.780464883e-07 wk1 = 1.492301901e-07 pk1 = -1.883406599e-13
+ k2 = -6.586573078e-02 lk2 = 1.056693295e-07 wk2 = -3.317794926e-08 pk2 = 1.677447726e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.328619896e+05 lvsat = -3.955383029e-01 wvsat = 1.975796604e-01 pvsat = -3.587930694e-7
+ ua = -1.106891114e-09 lua = -5.495446189e-16 wua = 4.089756758e-16 pua = 6.292675285e-23
+ ub = 2.583787673e-18 lub = 3.371850094e-25 wub = -7.234493320e-25 pub = 5.604985142e-31
+ uc = 1.153509676e-10 luc = 3.534849816e-17 wuc = -1.945799790e-16 puc = 1.262691162e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.554241413e-02 lu0 = -4.682656412e-09 wu0 = -7.287713461e-09 pu0 = 8.909308249e-15
+ a0 = 9.810135182e-01 la0 = 1.681865498e-06 wa0 = 1.610519426e-06 pa0 = -3.119869886e-12
+ keta = 3.313231538e-01 lketa = -1.317324293e-06 wketa = -2.433313664e-07 pketa = 9.674733464e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -1.073353111e+00 lags = 6.386582974e-06 wags = 1.130089584e-06 pags = -4.466332890e-12
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.214881825e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 5.065702825e-09 wvoff = 2.872873883e-08 pvoff = -5.081537924e-14
+ nfactor = {5.322684447e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.519801001e-06 wnfactor = 2.423799404e-06 pnfactor = -4.714206196e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -9.185185185e-07 wcit = 1.744779259e-11
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386811553e-01 letab = 2.730728394e-07 wetab = 2.699468120e-11 petab = -1.073295027e-16
+ dsub = 8.410209171e-01 ldsub = -1.117325115e-06 wdsub = -2.000073164e-07 pdsub = 7.952190897e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.754186890e-01 lpclm = -2.998609364e-07 wpclm = -1.750344782e-07 ppclm = 6.959283337e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 7.840045856e-03 lpdiblc2 = -8.523204859e-09 wpdiblc2 = -7.030552144e-09 ppdiblc2 = 3.985173222e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.052861340e-05 lalpha0 = 5.005988890e-10 walpha0 = 8.079180259e-11 palpha0 = -2.808357176e-16
+ alpha1 = 0.0
+ beta0 = 1.384674463e+01 lbeta0 = 1.571228195e-05 wbeta0 = 9.421900382e-07 pbeta0 = -3.779218461e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.714177674e-01 lkt1 = 7.070807688e-08 wkt1 = 3.922581063e-08 pkt1 = -1.813498494e-13
+ kt2 = -3.059006496e-02 lkt2 = -9.204118984e-09 wkt2 = -8.082129757e-09 pkt2 = 1.015723646e-14
+ at = 1.210867672e+06 lat = -2.323262024e+00 wat = -1.827614374e+00 pat = 3.655714141e-6
+ ute = -1.393860885e+00 lute = 1.507992271e-07 wute = 2.440075888e-07 pute = 1.425577048e-13
+ ua1 = 2.015173602e-09 lua1 = 8.481085314e-16 wua1 = -2.129800571e-16 pua1 = -8.361557683e-22
+ ub1 = -2.439966397e-18 lub1 = -1.534024486e-24 wub1 = 2.232591510e-24 pub1 = -2.371392589e-31
+ uc1 = -2.478492555e-10 luc1 = 2.804466520e-16 wuc1 = 6.120375845e-16 puc1 = -9.039268787e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.43 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.387426635e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.109271451e-09 wvth0 = -1.497097716e-08 pvth0 = 1.942114569e-14
+ k1 = 4.338163653e-01 lk1 = -1.901770380e-08 wk1 = 3.923539383e-08 pk1 = 2.900355780e-14
+ k2 = -9.446557747e-03 lk2 = -5.812135502e-09 wk2 = -2.203802108e-08 pk2 = -5.237463814e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.809722383e+03 lvsat = 7.408911645e-02 wvsat = 1.135434016e-02 pvsat = 9.178852168e-9
+ ua = -1.308796443e-09 lua = -1.505897834e-16 wua = 9.441221524e-16 pua = -9.944959277e-22
+ ub = 2.817887276e-18 lub = -1.253841006e-25 wub = -7.413920635e-25 pub = 5.959524545e-31
+ uc = 1.580311898e-10 luc = -4.898548689e-17 wuc = -1.594818452e-16 puc = 5.691695868e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.580643157e-02 lu0 = -5.204341672e-09 wu0 = 5.494252934e-10 pu0 = -6.576486073e-15
+ a0 = 2.022100541e+00 la0 = -3.752704044e-07 wa0 = 3.092695612e-07 pa0 = -5.486652154e-13
+ keta = -3.973934933e-01 lketa = 1.225833655e-07 wketa = 2.382557425e-07 pketa = 1.588129847e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.835185489e+00 lags = 6.394561276e-07 wags = -1.026024682e-06 pags = -2.059589072e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.205835450e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.278184295e-09 wvoff = 2.716023694e-09 pvoff = 5.844452425e-16
+ nfactor = {8.530746986e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.859038833e-07 wnfactor = -1.908826884e-07 pnfactor = 4.522748856e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.694696667e-06 lcit = 1.141343921e-11 wcit = 3.447596577e-11 pcit = -3.364681880e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.960189626e-04 leta0 = 7.866330862e-12 weta0 = 1.101041678e-10 peta0 = -2.175603303e-16
+ etab = -4.918386561e-04 letab = 1.765917598e-11 wetab = -5.685009550e-11 petab = 5.834358379e-17
+ dsub = -4.674238962e-01 ldsub = 1.468096414e-06 wdsub = 1.123839262e-06 pdsub = -1.820635556e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.972782026e-01 lpclm = -3.430542424e-07 wpclm = -6.500979299e-08 ppclm = 4.785250569e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -4.249112654e-03 lpdiblc2 = 1.536436790e-08 wpdiblc2 = 2.097045797e-08 ppdiblc2 = -1.547686371e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.753434331e-04 lalpha0 = -2.223459813e-10 walpha0 = -1.204783304e-10 palpha0 = 1.168640018e-16
+ alpha1 = 0.0
+ beta0 = 2.271538963e+01 lbeta0 = -1.811717144e-06 wbeta0 = -1.783241126e-06 pbeta0 = 1.606097248e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.118014028e-01 lkt1 = -4.709087883e-08 wkt1 = -8.906115459e-08 pkt1 = 7.213877950e-14
+ kt2 = -5.124450336e-02 lkt2 = 3.160801858e-08 wkt2 = 2.017029381e-10 pkt2 = -6.211202750e-15
+ at = -4.285565109e+03 lat = 7.782001402e-02 wat = 3.960351870e-02 pat = -3.381505289e-8
+ ute = -1.508226546e+00 lute = 3.767800553e-07 wute = 5.790689957e-07 pute = -5.195068822e-13
+ ua1 = 1.382030307e-09 lua1 = 2.099168025e-15 wua1 = 1.140573072e-15 pua1 = -3.510709073e-21
+ ub1 = -1.827962019e-18 lub1 = -2.743314536e-24 wub1 = -3.691072323e-25 pub1 = 4.903687371e-30
+ uc1 = -7.983394413e-11 luc1 = -5.154320262e-17 wuc1 = 1.764676197e-16 puc1 = -4.326240667e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.44 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.427000038e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -6.971437699e-09 wvth0 = 6.699992964e-09 pvth0 = -1.728637604e-15
+ k1 = 4.458492289e-01 lk1 = -3.076117699e-08 wk1 = -4.854736623e-09 pk1 = 7.203332062e-14
+ k2 = -2.111234221e-02 lk2 = 5.573086843e-09 wk2 = -3.221914327e-09 pk2 = -2.360104320e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -1.930420324e+04 lvsat = 8.823500504e-02 wvsat = 3.214521158e-02 pvsat = -1.111199879e-8
+ ua = -2.322253647e-09 lua = 8.384937747e-16 wua = 1.810003609e-15 pua = -1.839552935e-21
+ ub = 3.672431807e-18 lub = -9.593768357e-25 wub = -1.772243561e-24 pub = 1.602011973e-30
+ uc = 1.739231150e-10 luc = -6.449521130e-17 wuc = -2.253642919e-16 puc = 1.212149326e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.586542154e-02 lu0 = 4.497587064e-09 wu0 = 7.307878148e-09 pu0 = -1.317239814e-14
+ a0 = 5.436060460e-01 la0 = 1.067666298e-06 wa0 = 2.257639409e-06 pa0 = -2.450176768e-12
+ keta = -5.053476732e-01 lketa = 2.279412473e-07 wketa = 4.566115679e-07 pketa = -1.972230693e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.436316423e+00 lags = -9.231676077e-07 wags = -4.824758967e-07 pags = -7.364353440e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.361905003e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.850979239e-08 wvoff = 4.530212557e-08 pvoff = -4.097746089e-14
+ nfactor = {8.855102774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.542483801e-07 wnfactor = 1.078443408e-06 pnfactor = -7.865239178e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 4.016844969e-03 leta0 = -3.428283810e-09 weta0 = -9.189356519e-09 peta0 = 8.858248327e-15
+ etab = -8.589439784e-04 letab = 3.759356153e-10 wetab = 9.078293831e-11 petab = -8.573887555e-17
+ dsub = 1.071928124e+00 ldsub = -3.423419066e-08 wdsub = -1.447649257e-06 pdsub = 6.890086641e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.512607821e-01 lpclm = 2.898873798e-07 wpclm = 7.281809788e-07 ppclm = -2.955894768e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 8.020941525e-03 lpdiblc2 = 3.389408521e-09 wpdiblc2 = 2.183834556e-08 ppdiblc2 = -1.632387861e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.352635408e-05 lalpha0 = 2.341489699e-11 walpha0 = -1.050468430e-10 palpha0 = 1.018036417e-16
+ alpha1 = 0.0
+ beta0 = 1.871845064e+01 lbeta0 = 2.089095470e-06 wbeta0 = -2.058391123e-06 pbeta0 = 1.874629888e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.755042347e-01 lkt1 = 1.507989996e-08 wkt1 = 1.129613363e-08 pkt1 = -2.580491594e-14
+ kt2 = -2.533845432e-02 lkt2 = 6.325010018e-09 wkt2 = 2.409490291e-08 pkt2 = -2.952977126e-14
+ at = 8.961427625e+04 lat = -1.382153615e-02 wat = -2.200050967e-02 pat = 2.630739860e-8
+ ute = -2.567642377e-01 lute = -8.445845847e-07 wute = -1.280927704e-06 pute = 1.295756897e-12
+ ua1 = 7.928871160e-09 lua1 = -4.290221305e-15 wua1 = -8.668015787e-15 pua1 = 6.061983223e-21
+ ub1 = -1.037333244e-17 lub1 = 5.596539723e-24 wub1 = 1.315966389e-23 pub1 = -8.299716807e-30
+ uc1 = -2.721042218e-10 luc1 = 1.361029749e-16 wuc1 = 2.968062796e-16 puc1 = -1.607069218e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.45 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.957984717e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.224365347e-08 wvth0 = -3.237390248e-10 pvth0 = 1.614307636e-15
+ k1 = 2.033435329e-01 lk1 = 8.465940904e-08 wk1 = 2.464172108e-07 pk1 = -4.755956275e-14
+ k2 = 5.016850393e-02 lk2 = -2.835303188e-08 wk2 = -9.903252526e-08 pk2 = 2.200001707e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.551563070e+05 lvsat = 5.200525174e-03 wvsat = 5.888276663e-02 pvsat = -2.383773811e-8
+ ua = 6.913796266e-10 lua = -5.958449818e-16 wua = -3.565762175e-15 pua = 7.190427899e-22
+ ub = 6.281798160e-19 lub = 4.895348993e-25 wub = 3.183262384e-24 pub = -7.565610809e-31
+ uc = 2.412569375e-11 luc = 6.800871330e-18 wuc = 7.371553284e-17 puc = -2.113211000e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.641312989e-02 lu0 = -5.282094728e-09 wu0 = -3.134728962e-08 pu0 = 5.225528964e-15
+ a0 = 3.976389470e+00 la0 = -5.661669730e-07 wa0 = -5.566202298e-06 pa0 = 1.273580692e-12
+ keta = -1.372235289e-02 lketa = -6.047823863e-09 wketa = 6.107735398e-08 pketa = -8.968560223e-15
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.849388776e+00 lags = -6.438193940e-07 wags = -3.864278988e-06 pags = 8.731338374e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.616877341e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -5.298048535e-09 wvoff = -7.476383756e-08 pvoff = 1.616793427e-14
+ nfactor = {2.954877863e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.306671224e-07 wnfactor = -1.385195526e-06 pnfactor = 3.860450325e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.034915704e-05 lcit = -2.545931292e-12 wcit = -1.576931495e-11 pcit = 7.505405448e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.919342104e-02 leta0 = 7.618642295e-09 weta0 = 3.477250968e-08 peta0 = -1.206540189e-14
+ etab = 2.738833180e-02 letab = -1.306835529e-08 wetab = -3.171597865e-08 petab = 1.505268930e-14
+ dsub = 1.756176225e+00 ldsub = -3.599020741e-07 wdsub = -2.686674326e-07 pdsub = 1.278722645e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.735387542e-01 lpclm = -5.508095956e-08 wpclm = -4.156632718e-07 ppclm = 2.488231943e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 8.259700170e-03 lpdiblc2 = 3.275771344e-09 wpdiblc2 = -8.637899337e-09 ppdiblc2 = -1.818709848e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.313527983e-03 lalpha0 = 1.135735909e-09 walpha0 = 2.080880250e-09 palpha0 = -9.385883582e-16
+ alpha1 = 0.0
+ beta0 = 1.587825466e+01 lbeta0 = 3.440886743e-06 wbeta0 = 5.276494974e-06 pbeta0 = -1.616409150e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.194818870e-01 lkt1 = -1.158393640e-08 wkt1 = -8.102023469e-08 pkt1 = 1.813305956e-14
+ kt2 = -1.247697135e-02 lkt2 = 2.035871961e-10 wkt2 = -5.360157090e-08 pkt2 = 7.449865448e-15
+ at = 6.087928044e+04 lat = -1.451148972e-04 wat = 7.359507879e-02 pat = -1.919132173e-8
+ ute = -1.619708861e+00 lute = -1.958910911e-07 wute = 6.262630413e-07 pute = 3.880294617e-13
+ ua1 = -8.740234288e-10 lua1 = -1.004836256e-16 wua1 = 4.197274343e-15 pua1 = -6.125161386e-23
+ ub1 = 1.594766595e-18 lub1 = -9.967701081e-26 wub1 = -5.238539439e-24 pub1 = 4.569080685e-31
+ uc1 = 9.361701639e-11 luc1 = -3.796204845e-17 wuc1 = -1.956485676e-16 puc1 = 7.367696269e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.46 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.042741516e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -3.415873336e-08 wvth0 = 1.883619221e-07 pvth0 = -4.101921749e-14
+ k1 = 4.231890419e-01 lk1 = 3.498531627e-08 wk1 = -1.787441287e-07 pk1 = 4.850564191e-14
+ k2 = -3.326318561e-02 lk2 = -9.501641625e-09 wk2 = 5.693075422e-08 pk2 = -1.323988593e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.009298497e+05 lvsat = -5.142006783e-03 wvsat = -1.233074270e-01 pvsat = 1.732813614e-8
+ ua = -1.320720833e-09 lua = -1.412108828e-16 wua = -1.107189159e-15 pua = 1.635282169e-22
+ ub = 2.606970466e-18 lub = 4.242715188e-26 wub = 9.498074711e-25 pub = -2.519119434e-31
+ uc = 6.670078480e-11 luc = -2.818970493e-18 wuc = -6.858026216e-19 puc = -4.321128252e-24
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.271971214e-02 lu0 = -2.188066985e-09 wu0 = -1.109413382e-08 pu0 = 6.493284110e-16
+ a0 = 4.747117541e+00 la0 = -7.403129805e-07 wa0 = 2.271040419e-07 pa0 = -3.541687534e-14
+ keta = 1.378862962e-01 lketa = -4.030379812e-08 wketa = 6.151524964e-09 pketa = 3.441930842e-15
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.667043698e+00 lags = 6.026185235e-07 wags = 3.653891799e-07 pags = -8.255968521e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.362495478e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 6.017702427e-09 wvoff = -4.481114241e-08 pvoff = 9.400122796e-15
+ nfactor = {1.522449504e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.929900653e-07 wnfactor = -5.663973127e-07 pnfactor = 2.010375763e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.410413228e-05 lcit = 2.979289428e-12 wcit = 5.631898195e-11 pcit = -8.782945235e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.470592107e-01 leta0 = 3.650991748e-08 weta0 = -1.495964464e-08 peta0 = -8.284216229e-16
+ etab = -7.892538262e-02 letab = 1.095322848e-08 wetab = 1.528774307e-07 petab = -2.665619153e-14
+ dsub = -2.109379238e-01 ldsub = 8.456736774e-08 wdsub = 9.325907543e-07 pdsub = -1.435520228e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 3.304620937e-02 lpclm = 2.185333095e-08 wpclm = 1.962662683e-06 ppclm = -2.885595553e-13
+ pdiblc1 = -9.545380289e-01 lpdiblc1 = 3.037983676e-07 wpdiblc1 = -2.309881556e-08 ppdiblc1 = 5.219177376e-15
+ pdiblc2 = 5.153298225e-02 lpdiblc2 = -6.501826742e-09 wpdiblc2 = -7.010385725e-08 ppdiblc2 = 1.206952334e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.351877991e-03 lalpha0 = -1.048162571e-09 walpha0 = -6.127014504e-09 palpha0 = 9.159854614e-16
+ alpha1 = 0.0
+ beta0 = 3.577380792e+01 lbeta0 = -1.054513515e-06 wbeta0 = -3.677006707e-06 pbeta0 = 4.066345551e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.045905124e-01 lkt1 = -1.494864250e-08 wkt1 = 1.081591155e-08 pkt1 = -2.617317680e-15
+ kt2 = 1.386596703e-02 lkt2 = -5.748599731e-09 wkt2 = -7.420254313e-08 pkt2 = 1.210465512e-14
+ at = 4.696992662e+04 lat = 2.997703600e-03 wat = -6.453240070e-02 pat = 1.201858226e-8
+ ute = -4.280884613e+00 lute = 4.054015700e-07 wute = 7.843083371e-06 pute = -1.242611092e-12
+ ua1 = -4.764604935e-09 lua1 = 7.785932657e-16 wua1 = 1.433403599e-14 pua1 = -2.351652909e-21
+ ub1 = 3.768904403e-18 lub1 = -5.909234485e-25 wub1 = -1.203122565e-23 pub1 = 1.991715517e-30
+ uc1 = -1.828714253e-10 luc1 = 2.451051494e-17 wuc1 = 2.914556219e-16 puc1 = -3.638422893e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.47 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.65e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.547334207e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -4.202785638e-08 wvth0 = -5.770991457e-07 pvth0 = 7.835443603e-14
+ k1 = 6.445692952e-01 lk1 = 4.610657745e-10 wk1 = 6.876831679e-07 pk1 = -8.661369500e-14
+ k2 = -1.274477187e-01 lk2 = 5.186436309e-09 wk2 = -1.694110344e-07 pk2 = 2.205811602e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.803657937e+05 lvsat = -1.935042249e-03 wvsat = -7.848529550e-02 pvsat = 1.033812473e-8
+ ua = -1.607991728e-09 lua = -9.641098684e-17 wua = -2.512115080e-16 pua = 3.003850219e-23
+ ub = 3.756687818e-18 lub = -1.368712691e-25 wub = -2.601168913e-24 pub = 3.018628238e-31
+ uc = 1.360461490e-10 luc = -1.363338004e-17 wuc = -1.476026390e-16 puc = 1.859055239e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.785910730e-02 lu0 = -2.989555662e-09 wu0 = -2.965822690e-08 pu0 = 3.544398727e-15
+ a0 = 0.0
+ keta = 1.118741745e-01 lketa = -3.624720774e-08 wketa = 1.467087053e-07 pketa = -1.847796144e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 9.861009617e-01 lags = 3.291061387e-08 wags = -8.525747532e-07 pags = 1.073817902e-13
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.618938198e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.001692666e-08 wvoff = 8.039417125e-08 pvoff = -1.012564587e-14
+ nfactor = {1.916882308e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 4.005222859e-07 wnfactor = 2.414960298e-06 pnfactor = -2.639051431e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.599166667e-05 lcit = 3.273650417e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.202815303e-01 leta0 = -5.181871083e-09 weta0 = -1.053792735e-07 peta0 = 1.327251949e-14
+ etab = -4.517283131e-02 letab = 5.689518104e-09 wetab = -9.383187403e-08 petab = 1.181812453e-14
+ dsub = 6.308199508e-01 ldsub = -4.670477281e-08 wdsub = 6.285017821e-08 pdsub = -7.915979946e-15
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.948675935e-01 lpclm = -3.382713899e-09 wpclm = 5.839230065e-07 ppclm = -7.354510267e-14
+ pdiblc1 = 9.662720674e-01 lpdiblc1 = 4.248033112e-09 wpdiblc1 = 5.389723631e-08 ppdiblc1 = -6.788356913e-15
+ pdiblc2 = 2.666624417e-02 lpdiblc2 = -2.623858938e-09 wpdiblc2 = 3.789422680e-08 ppdiblc2 = -4.772777865e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.875110871e-03 lalpha0 = -1.940607386e-10 walpha0 = -1.317415016e-09 palpha0 = 1.659284213e-16
+ alpha1 = 0.0
+ beta0 = 3.341427165e+01 lbeta0 = -6.865438332e-07 wbeta0 = -5.559821364e-06 pbeta0 = 7.002595008e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -6.821869689e-02 lkt1 = -3.621582713e-08 wkt1 = -3.101920910e-08 pkt1 = 3.906869387e-15
+ kt2 = -7.062948907e-02 lkt2 = 7.428466649e-09 wkt2 = 1.775895071e-08 pkt2 = -2.236739842e-15
+ at = -2.153146649e+04 lat = 1.368049585e-02 wat = 6.515847901e-02 pat = -8.206710431e-9
+ ute = -1.756571846e+00 lute = 1.173499403e-08 wute = -6.494080035e-07 pute = 8.179293804e-14
+ ua1 = 5.428011876e-10 lua1 = -4.909671907e-17 wua1 = -3.875333191e-15 pua1 = 4.880982154e-22
+ ub1 = 2.282776272e-19 lub1 = -3.876270290e-26 wub1 = 3.848195918e-24 pub1 = -4.846802759e-31
+ uc1 = 3.099879242e-11 luc1 = -8.842545505e-18 wuc1 = 3.022758438e-16 puc1 = -3.807164252e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.48 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.49 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.50 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.120860594e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.320442463e-8
+ k1 = 6.076841567e-01 lk1 = -2.959067260e-7
+ k2 = -8.662790178e-02 lk2 = 1.161664992e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.565038297e+05 lvsat = -6.200646292e-1
+ ua = -8.509614041e-10 lua = -5.101661753e-16
+ ub = 2.131065938e-18 lub = 6.879350183e-25
+ uc = -6.413725184e-12 luc = 1.143654670e-16 puc = 2.350988702e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.098189256e-02 lu0 = 8.926303521e-10
+ a0 = 1.988847952e+00 la0 = -2.704936295e-7
+ keta = 1.790507093e-01 lketa = -7.118966674e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.661631337e-01 lags = 3.591631228e-06 pags = 8.077935669e-28
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.035102483e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.673365840e-8
+ nfactor = {2.049039036e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.430265455e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 7.158598930e-01 ldsub = -6.196911417e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.658852232e-01 lpclm = 1.356386466e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.440451272e-03 lpdiblc2 = 1.641530091e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.997053919e-05 lalpha0 = 3.248568880e-10
+ alpha1 = 0.0
+ beta0 = 1.443635041e+01 lbeta0 = 1.334731420e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.468709522e-01 lkt1 = -4.277743590e-8
+ kt2 = -3.564771813e-02 lkt2 = -2.847900921e-9
+ at = 6.717907755e+04 lat = -3.558108488e-2
+ ute = -1.241165272e+00 lute = 2.400093052e-7
+ ua1 = 1.881894467e-09 lua1 = 3.248571119e-16
+ ub1 = -1.042850307e-18 lub1 = -1.682422020e-24
+ uc1 = 1.351529876e-10 luc1 = -2.852147239e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.51 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.293740921e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 9.044136365e-9
+ k1 = 4.583691775e-01 lk1 = -8.677927811e-10
+ k2 = -2.323755968e-02 lk2 = -9.089647275e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.295621900e+03 lvsat = 7.983307901e-2
+ ua = -7.179815791e-10 lua = -7.729276606e-16
+ ub = 2.353937298e-18 lub = 2.475523540e-25
+ uc = 5.823028540e-11 luc = -1.336786569e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.615025215e-02 lu0 = -9.319789778e-9
+ a0 = 2.215635936e+00 la0 = -7.186153452e-7
+ keta = -2.482972840e-01 lketa = 1.325215998e-07 wketa = 1.058791184e-22
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.193117478e+00 lags = 5.105707038e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.188839056e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.643919741e-9
+ nfactor = {7.336237045e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.168929469e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.487975000e-05 lcit = -9.642142012e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.649201940e-04 leta0 = -1.282790573e-10
+ etab = -5.274144355e-04 letab = 5.416955383e-11
+ dsub = 2.358547406e-01 ldsub = 3.287750393e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.565962295e-01 lpclm = -4.360176618e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.873827250e-03 lpdiblc2 = 5.679221645e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.999502351e-04 lalpha0 = -1.492145659e-10
+ alpha1 = 0.0
+ beta0 = 2.159946903e+01 lbeta0 = -8.066500302e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.675342905e-01 lkt1 = -1.947712687e-9
+ kt2 = -5.111828125e-02 lkt2 = 2.772115829e-8
+ at = 2.049761305e+04 lat = 5.665915489e-2
+ ute = -1.145855460e+00 lute = 5.168188119e-8
+ ua1 = 2.095780665e-09 lua1 = -9.777132001e-17
+ ub1 = -2.058942765e-18 lub1 = 3.253258715e-25
+ uc1 = 3.059635606e-11 luc1 = -7.861604784e-17 wuc1 = 6.162975822e-33 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.52 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.468927403e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -8.053188390e-9
+ k1 = 4.428112210e-01 lk1 = 1.431599487e-8
+ k2 = -2.312855893e-02 lk2 = -9.196026549e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.116988700e+02 lvsat = 8.128131369e-2
+ ua = -1.189585556e-09 lua = -3.126657592e-16
+ ub = 2.563393283e-18 lub = 4.313378596e-26
+ uc = 3.289414631e-11 luc = 1.135893926e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.043856181e-02 lu0 = -3.745465588e-9
+ a0 = 1.956396665e+00 la0 = -4.656107786e-7
+ keta = -2.196082690e-01 lketa = 1.045225556e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.134391582e+00 lags = -1.384015758e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.078412353e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -7.133174371e-9
+ nfactor = {1.560380996e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.620556907e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.733691026e-03 leta0 = 2.115050563e-09 weta0 = 4.135903063e-25 peta0 = 1.972152263e-31
+ etab = -8.021336290e-04 letab = 3.222817507e-10
+ dsub = 1.660149467e-01 ldsub = 3.969351861e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044219330e-01 lpclm = 1.049127385e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.168699006e-02 lpdiblc2 = -6.825784599e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.221009338e-05 lalpha0 = 8.712180668e-11 palpha0 = 1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.743034605e+01 lbeta0 = 3.262205538e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.684353150e-01 lkt1 = -1.068357826e-9
+ kt2 = -1.026029230e-02 lkt2 = -1.215419603e-8
+ at = 7.584674830e+04 lat = 2.641166347e-3
+ ute = -1.058346030e+00 lute = -3.372294702e-8
+ ua1 = 2.504580930e-09 lua1 = -4.967399386e-16
+ ub1 = -2.138248650e-18 lub1 = 4.027244500e-25
+ uc1 = -8.636812690e-11 luc1 = 3.553543930e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.53 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955958815e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.123344844e-8
+ k1 = 3.575470440e-01 lk1 = 5.489747991e-8
+ k2 = -1.180429035e-02 lk2 = -1.458581218e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.920040959e+05 lvsat = -9.716707688e-3
+ ua = -1.540010971e-09 lua = -1.458807828e-16
+ ub = 2.620208842e-18 lub = 1.609242065e-26
+ uc = 7.025556412e-11 luc = -6.423227544e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.679655316e-02 lu0 = -2.012051571e-9
+ a0 = 4.931589960e-01 la0 = 2.308171899e-7
+ keta = 2.449876974e-02 lketa = -1.166018946e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.311916620e-01 lags = -9.742775603e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.329546542e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.819557388e-9
+ nfactor = {2.088047121e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.109129981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.810000000e-07 lcit = 2.150818050e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.566597539e-03 leta0 = 6.832822021e-11
+ etab = 7.541036029e-03 letab = -3.648649848e-09 wetab = 1.344168495e-24 petab = 4.683861625e-31
+ dsub = 1.588048920e+00 ldsub = -2.798818835e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.134240660e-01 lpclm = 1.006281733e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.854256280e-03 lpdiblc2 = 2.137655044e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.011350105e-03 lalpha0 = 5.483839952e-10
+ alpha1 = 0.0
+ beta0 = 1.918019144e+01 lbeta0 = 2.429366624e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701829100e-01 lkt1 = -2.365899855e-10
+ kt2 = -4.601988180e-02 lkt2 = 4.865580593e-9
+ at = 1.069337728e+05 lat = -1.215470296e-2
+ ute = -1.227804580e+00 lute = 4.693084985e-8
+ ua1 = 1.752556260e-09 lua1 = -1.388137969e-16
+ ub1 = -1.683418286e-18 lub1 = 1.862479382e-25 wub1 = 7.346839693e-40
+ uc1 = -2.881638008e-11 luc1 = 8.143685399e-18 wuc1 = -6.162975822e-33 puc1 = -1.469367939e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.54 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.221476949e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.982783066e-8
+ k1 = 3.113341429e-01 lk1 = 6.533928492e-8
+ k2 = 2.363068596e-03 lk2 = -1.778692694e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.237662533e+05 lvsat = 5.701632855e-3
+ ua = -2.013580132e-09 lua = -3.887783096e-17
+ ub = 3.201343101e-18 lub = -1.152148652e-25
+ uc = 6.627162171e-11 luc = -5.523055757e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.577720036e-02 lu0 = -1.781728806e-9
+ a0 = 4.889235214e+00 la0 = -7.624762317e-7
+ keta = 1.417358112e-01 lketa = -3.814989897e-08 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.438389643e+00 lags = 5.509541398e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.642915643e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.190013221e-8
+ nfactor = {1.168008132e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.187958077e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.113928571e-05 lcit = -2.516921607e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.564206905e-01 leta0 = 3.599150595e-08 weta0 = -3.308722450e-24 peta0 = 1.577721810e-30
+ etab = 1.674259653e-02 letab = -5.727742443e-9
+ dsub = 3.726607961e-01 ldsub = -5.264936889e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.261245636e+00 lpclm = -1.587221104e-7
+ pdiblc1 = -9.689928571e-01 lpdiblc1 = 3.070644361e-7
+ pdiblc2 = 7.663234286e-03 lpdiblc2 = 1.051066463e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.517701205e-03 lalpha0 = -4.749551482e-10
+ alpha1 = 0.0
+ beta0 = 3.347280247e+01 lbeta0 = -8.000488374e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.978221071e-01 lkt1 = -1.658651339e-8
+ kt2 = -3.256866571e-02 lkt2 = 1.826278318e-9
+ at = 6.586697143e+03 lat = 1.051871878e-2
+ ute = 6.271775714e-01 lute = -3.722023673e-7
+ ua1 = 4.205380043e-09 lua1 = -6.930293307e-16 pua1 = -1.880790961e-37
+ ub1 = -3.760022786e-18 lub1 = 6.554567249e-25
+ uc1 = -4.836768571e-13 luc1 = 1.741911106e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.55 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1e-06 wmax = 1.65e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.199425423e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -1.269893712e-08 wvth0 = -2.019033219e-07 pvth0 = 3.148682306e-14
+ k1 = 1.162898258e+00 lk1 = -6.746213876e-08 wk1 = -1.406065139e-07 pk1 = 2.192758585e-14
+ k2 = -2.675054486e-01 lk2 = 2.429906832e-08 wk2 = 5.440121798e-08 pk2 = -8.483869943e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 7.842422391e+04 lvsat = 1.277272234e-02 wvsat = 8.441733297e-02 pvsat = -1.316488308e-8
+ ua = -9.557611658e-11 lua = -3.379905572e-16 wua = -2.668051655e-15 pua = 4.160826556e-22
+ ub = 1.344944324e-18 lub = 1.742905241e-25 wub = 1.252797190e-24 pub = -1.953737218e-31
+ uc = -6.738595665e-11 luc = 1.532084359e-17 wuc = 1.774818658e-16 puc = -2.767829697e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 4.308038042e-02 lu0 = -4.480159737e-09 wu0 = -3.800182135e-08 pu0 = 5.926384040e-15
+ a0 = 0.0
+ keta = 1.280836202e+00 lketa = -2.157926049e-07 wketa = -1.721292615e-06 pketa = 2.684355833e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.427778610e-01 lags = 1.016360676e-07 wags = 1.565556175e-08 pags = -2.441484855e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.986804670e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.285808158e-08 wvoff = 2.989792333e-07 pvoff = -4.662581144e-14
+ nfactor = {3.513481879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 4.461539260e-07 wnfactor = 2.159823686e-06 pnfactor = -3.368245039e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.599166667e-05 lcit = 3.273650417e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.362264692e-01 leta0 = 3.284221713e-08 weta0 = 3.045205096e-07 peta0 = -4.748997348e-14
+ etab = -1.754397557e-01 letab = 2.424309539e-08 wetab = 1.143346712e-07 petab = -1.783049197e-14
+ dsub = 6.701504754e-01 ldsub = -5.165845237e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.554362767e+00 lpclm = -2.044337270e-07 wpclm = -1.588550281e-06 ppclm = 2.477344163e-13
+ pdiblc1 = 6.937249699e-01 lpdiblc1 = 4.776359095e-08 wpdiblc1 = 4.894274982e-07 ppdiblc1 = -7.632621834e-14
+ pdiblc2 = 6.081967645e-02 lpdiblc2 = -7.238680692e-09 wpdiblc2 = -1.668295799e-08 ppdiblc2 = 2.601707298e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.411199537e-04 lalpha0 = 5.162269786e-11 walpha0 = 1.453502470e-09 palpha0 = -2.266737102e-16
+ alpha1 = 0.0
+ beta0 = 2.333846338e+01 lbeta0 = 7.804013446e-07 wbeta0 = 1.054132025e-05 pbeta0 = -1.643918893e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.961051924e-01 lkt1 = -9.361447576e-08 wkt1 = -6.132087842e-07 pkt1 = 9.562990990e-14
+ kt2 = -3.670706487e-02 lkt2 = 2.471661666e-09 wkt2 = -3.644908317e-08 pkt2 = 5.684234520e-15
+ at = -6.217541132e+04 lat = 2.124216960e-02 wat = 1.301075028e-01 pat = -2.029026507e-8
+ ute = -2.107239553e+00 lute = 5.422998334e-08 wute = -8.904100744e-08 pute = 1.388594511e-14
+ ua1 = -3.498691419e-09 lua1 = 5.084206137e-16 wua1 = 2.582971994e-15 pua1 = -4.028144824e-22
+ ub1 = 5.418229913e-18 lub1 = -7.758917834e-25 wub1 = -4.445347835e-24 pub1 = 6.932519948e-31
+ uc1 = 3.799707541e-10 luc1 = -5.758995740e-17 wuc1 = -2.553813510e-16 puc1 = 3.982672169e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.56 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.57 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.58 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.120860594e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.320442463e-8
+ k1 = 6.076841567e-01 lk1 = -2.959067260e-7
+ k2 = -8.662790178e-02 lk2 = 1.161664992e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.565038297e+05 lvsat = -6.200646292e-1
+ ua = -8.509614041e-10 lua = -5.101661753e-16
+ ub = 2.131065938e-18 lub = 6.879350183e-25
+ uc = -6.413725184e-12 luc = 1.143654670e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.098189256e-02 lu0 = 8.926303521e-10
+ a0 = 1.988847952e+00 la0 = -2.704936295e-7
+ keta = 1.790507092e-01 lketa = -7.118966674e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.661631336e-01 lags = 3.591631228e-06 pags = -1.615587134e-27
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.035102483e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.673365840e-8
+ nfactor = {2.049039036e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.430265455e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 7.158598930e-01 ldsub = -6.196911417e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.658852232e-01 lpclm = 1.356386466e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.440451272e-03 lpdiblc2 = 1.641530091e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.997053919e-05 lalpha0 = 3.248568880e-10
+ alpha1 = 0.0
+ beta0 = 1.443635041e+01 lbeta0 = 1.334731420e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.468709523e-01 lkt1 = -4.277743590e-8
+ kt2 = -3.564771813e-02 lkt2 = -2.847900921e-9
+ at = 6.717907755e+04 lat = -3.558108488e-2
+ ute = -1.241165272e+00 lute = 2.400093052e-7
+ ua1 = 1.881894468e-09 lua1 = 3.248571119e-16
+ ub1 = -1.042850307e-18 lub1 = -1.682422020e-24
+ uc1 = 1.351529876e-10 luc1 = -2.852147239e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.59 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.293740921e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 9.044136365e-9
+ k1 = 4.583691775e-01 lk1 = -8.677927811e-10
+ k2 = -2.323755967e-02 lk2 = -9.089647275e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.295621900e+03 lvsat = 7.983307901e-2
+ ua = -7.179815791e-10 lua = -7.729276606e-16
+ ub = 2.353937298e-18 lub = 2.475523540e-25
+ uc = 5.823028540e-11 luc = -1.336786569e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.615025215e-02 lu0 = -9.319789778e-9
+ a0 = 2.215635936e+00 la0 = -7.186153452e-7
+ keta = -2.482972840e-01 lketa = 1.325215998e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.193117478e+00 lags = 5.105707038e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.188839056e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.643919741e-9
+ nfactor = {7.336237045e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.168929469e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.487975000e-05 lcit = -9.642142013e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.649201940e-04 leta0 = -1.282790573e-10
+ etab = -5.274144355e-04 letab = 5.416955383e-11
+ dsub = 2.358547406e-01 ldsub = 3.287750393e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.565962295e-01 lpclm = -4.360176618e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.873827250e-03 lpdiblc2 = 5.679221645e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.999502351e-04 lalpha0 = -1.492145659e-10
+ alpha1 = 0.0
+ beta0 = 2.159946903e+01 lbeta0 = -8.066500302e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.675342905e-01 lkt1 = -1.947712687e-9
+ kt2 = -5.111828125e-02 lkt2 = 2.772115829e-8
+ at = 2.049761305e+04 lat = 5.665915489e-2
+ ute = -1.145855460e+00 lute = 5.168188119e-8
+ ua1 = 2.095780665e-09 lua1 = -9.777132001e-17
+ ub1 = -2.058942765e-18 lub1 = 3.253258715e-25
+ uc1 = 3.059635605e-11 luc1 = -7.861604784e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.60 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.468927403e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -8.053188390e-9
+ k1 = 4.428112210e-01 lk1 = 1.431599487e-8
+ k2 = -2.312855893e-02 lk2 = -9.196026549e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.116988700e+02 lvsat = 8.128131369e-2
+ ua = -1.189585556e-09 lua = -3.126657592e-16
+ ub = 2.563393283e-18 lub = 4.313378596e-26
+ uc = 3.289414631e-11 luc = 1.135893926e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.043856181e-02 lu0 = -3.745465588e-9
+ a0 = 1.956396665e+00 la0 = -4.656107786e-7
+ keta = -2.196082690e-01 lketa = 1.045225556e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.134391582e+00 lags = -1.384015758e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.078412353e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -7.133174371e-9
+ nfactor = {1.560380996e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.620556907e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.733691026e-03 leta0 = 2.115050563e-09 peta0 = -3.944304526e-31
+ etab = -8.021336290e-04 letab = 3.222817507e-10
+ dsub = 1.660149467e-01 ldsub = 3.969351861e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044219330e-01 lpclm = 1.049127385e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.168699006e-02 lpdiblc2 = -6.825784599e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.221009338e-05 lalpha0 = 8.712180668e-11 palpha0 = -2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.743034605e+01 lbeta0 = 3.262205538e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.684353150e-01 lkt1 = -1.068357826e-9
+ kt2 = -1.026029230e-02 lkt2 = -1.215419603e-8
+ at = 7.584674830e+04 lat = 2.641166347e-3
+ ute = -1.058346030e+00 lute = -3.372294702e-8
+ ua1 = 2.504580930e-09 lua1 = -4.967399386e-16
+ ub1 = -2.138248650e-18 lub1 = 4.027244500e-25
+ uc1 = -8.636812690e-11 luc1 = 3.553543930e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.61 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955958815e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.123344844e-8
+ k1 = 3.575470440e-01 lk1 = 5.489747991e-8
+ k2 = -1.180429035e-02 lk2 = -1.458581218e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.920040959e+05 lvsat = -9.716707688e-3
+ ua = -1.540010971e-09 lua = -1.458807828e-16
+ ub = 2.620208842e-18 lub = 1.609242065e-26
+ uc = 7.025556412e-11 luc = -6.423227544e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.679655316e-02 lu0 = -2.012051571e-09 wu0 = -2.646977960e-23
+ a0 = 4.931589960e-01 la0 = 2.308171899e-7
+ keta = 2.449876974e-02 lketa = -1.166018946e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.311916620e-01 lags = -9.742775603e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.329546542e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.819557388e-9
+ nfactor = {2.088047121e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.109129981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.810000000e-07 lcit = 2.150818050e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.566597539e-03 leta0 = 6.832822021e-11
+ etab = 7.541036029e-03 letab = -3.648649848e-09 wetab = 8.271806126e-25 petab = 7.888609052e-31
+ dsub = 1.588048920e+00 ldsub = -2.798818835e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.134240660e-01 lpclm = 1.006281733e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.854256280e-03 lpdiblc2 = 2.137655044e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.011350105e-03 lalpha0 = 5.483839952e-10 walpha0 = -4.135903063e-25 palpha0 = -9.860761315e-32
+ alpha1 = 0.0
+ beta0 = 1.918019144e+01 lbeta0 = 2.429366624e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701829100e-01 lkt1 = -2.365899855e-10
+ kt2 = -4.601988180e-02 lkt2 = 4.865580593e-9
+ at = 1.069337728e+05 lat = -1.215470296e-2
+ ute = -1.227804580e+00 lute = 4.693084985e-8
+ ua1 = 1.752556260e-09 lua1 = -1.388137969e-16
+ ub1 = -1.683418286e-18 lub1 = 1.862479382e-25
+ uc1 = -2.881638008e-11 luc1 = 8.143685399e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.62 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.221476949e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.982783066e-8
+ k1 = 3.113341429e-01 lk1 = 6.533928492e-8
+ k2 = 2.363068596e-03 lk2 = -1.778692694e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.237662533e+05 lvsat = 5.701632855e-3
+ ua = -2.013580132e-09 lua = -3.887783096e-17
+ ub = 3.201343101e-18 lub = -1.152148652e-25
+ uc = 6.627162171e-11 luc = -5.523055757e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.577720036e-02 lu0 = -1.781728806e-9
+ a0 = 4.889235214e+00 la0 = -7.624762317e-7
+ keta = 1.417358112e-01 lketa = -3.814989897e-08 pketa = -1.262177448e-29
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.438389643e+00 lags = 5.509541398e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.642915643e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.190013221e-8
+ nfactor = {1.168008132e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.187958077e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.113928571e-05 lcit = -2.516921607e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.564206905e-01 leta0 = 3.599150595e-08 peta0 = -7.888609052e-30
+ etab = 1.674259653e-02 letab = -5.727742443e-9
+ dsub = 3.726607961e-01 ldsub = -5.264936889e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.261245636e+00 lpclm = -1.587221104e-7
+ pdiblc1 = -9.689928571e-01 lpdiblc1 = 3.070644361e-7
+ pdiblc2 = 7.663234286e-03 lpdiblc2 = 1.051066463e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.517701205e-03 lalpha0 = -4.749551482e-10 walpha0 = -3.308722450e-24
+ alpha1 = 0.0
+ beta0 = 3.347280247e+01 lbeta0 = -8.000488374e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.978221071e-01 lkt1 = -1.658651339e-8
+ kt2 = -3.256866571e-02 lkt2 = 1.826278318e-9
+ at = 6.586697143e+03 lat = 1.051871878e-2
+ ute = 6.271775714e-01 lute = -3.722023673e-7
+ ua1 = 4.205380043e-09 lua1 = -6.930293307e-16
+ ub1 = -3.760022786e-18 lub1 = 6.554567249e-25 wub1 = 1.469367939e-39
+ uc1 = -4.836768571e-13 luc1 = 1.741911106e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.63 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.418104934e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 2.583495668e-07 wvth0 = 1.445765685e-06 pvth0 = -2.254671586e-13
+ k1 = 2.162141088e+00 lk1 = -2.232940581e-07 wk1 = -1.087888717e-06 pk1 = 1.696562454e-13
+ k2 = -4.030238912e-01 lk2 = 4.543316945e-08 wk2 = 1.828727016e-07 pk2 = -2.851899781e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.471012683e+05 lvsat = 2.062537256e-03 wvsat = 1.931149484e-02 pvsat = -3.011627621e-9
+ ua = -7.325503803e-09 lua = 7.895166655e-16 wua = 4.185919792e-15 pua = -6.527941915e-22
+ ub = 3.922161905e-18 lub = -2.276265576e-25 wub = -1.190405077e-24 pub = 1.856436717e-31
+ uc = 2.058877749e-11 luc = 1.601183799e-18 wuc = 9.408181780e-17 puc = -1.467205949e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -8.053582522e-02 lu0 = 1.479778753e-08 wu0 = 7.918634160e-08 pu0 = -1.234910997e-14
+ a0 = 0.0
+ keta = -2.764038217e+00 lketa = 4.150055607e-07 wketa = 2.113248334e-06 pketa = -3.295610777e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.034648292e-01 lags = 1.077669349e-07 wags = 5.292431595e-08 pags = -8.253547072e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {6.435719822e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.140861879e-07 wvoff = -5.942760885e-07 pvoff = 9.267735600e-14
+ nfactor = {1.349886398e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.604201162e-06 wnfactor = -1.030402129e-05 pnfactor = 1.606912120e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.599166667e-05 lcit = 3.273650417e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.046195544e-01 leta0 = 4.350811878e-08 weta0 = 3.693571545e-07 peta0 = -5.760124824e-14
+ etab = 1.438893247e-01 letab = -2.555627470e-08 wetab = -1.883892970e-07 petab = 2.937931087e-14
+ dsub = 6.709523213e-01 ldsub = -5.178350025e-08 wdsub = -7.601499898e-10 pdsub = 1.185453909e-16
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -1.287668283e-01 lpclm = 5.805033338e-08 wpclm = 7.056575460e-09 ppclm = -1.100472943e-15
+ pdiblc1 = 2.244242310e+00 lpdiblc1 = -1.940395882e-07 wpdiblc1 = -9.804629402e-07 ppdiblc1 = 1.529031955e-13
+ pdiblc2 = 2.750766875e-01 lpdiblc2 = -4.065206156e-08 wpdiblc2 = -2.197986045e-07 ppdiblc2 = 3.427759237e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -2.009620331e-03 lalpha0 = 3.870306452e-10 walpha0 = 3.492404260e-09 palpha0 = -5.446404443e-16
+ alpha1 = 0.0
+ beta0 = -9.551680915e+01 lbeta0 = 1.931588110e-05 wbeta0 = 1.232161186e-04 pbeta0 = -1.921555370e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -8.511178750e-01 lkt1 = 8.529496161e-08 wkt1 = 4.743586837e-07 pkt1 = -7.397623672e-14
+ kt2 = -3.143053049e-01 lkt2 = 4.576310720e-08 wkt2 = 2.267140484e-07 pkt2 = -3.535605585e-14
+ at = 1.509939690e+05 lat = -1.200159527e-02 wat = -7.197706969e-02 pat = 1.122482402e-8
+ ute = -3.642337046e+00 lute = 2.936284373e-07 wute = 1.366231415e-06 pute = -2.130637892e-13
+ ua1 = -3.178334752e-09 lua1 = 4.584609915e-16 wua1 = 2.279273874e-15 pua1 = -3.554527606e-22
+ ub1 = 1.790417750e-19 lub1 = 4.115960669e-26 wub1 = 5.214025201e-25 pub1 = -8.131272301e-32
+ uc1 = 7.747817220e-10 luc1 = -1.191607279e-16 wuc1 = -6.296621486e-16 puc1 = 9.819581208e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.64 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.65 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.66 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.120860594e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.320442463e-8
+ k1 = 6.076841567e-01 lk1 = -2.959067260e-7
+ k2 = -8.662790178e-02 lk2 = 1.161664992e-7
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.565038297e+05 lvsat = -6.200646292e-1
+ ua = -8.509614041e-10 lua = -5.101661753e-16
+ ub = 2.131065938e-18 lub = 6.879350183e-25
+ uc = -6.413725184e-12 luc = 1.143654670e-16 puc = 2.350988702e-38
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.098189256e-02 lu0 = 8.926303521e-10
+ a0 = 1.988847952e+00 la0 = -2.704936295e-7
+ keta = 1.790507092e-01 lketa = -7.118966674e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.661631337e-01 lags = 3.591631228e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.035102483e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.673365840e-8
+ nfactor = {2.049039036e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.430265455e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 7.158598930e-01 ldsub = -6.196911417e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.658852233e-01 lpclm = 1.356386466e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.440451272e-03 lpdiblc2 = 1.641530091e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.997053919e-05 lalpha0 = 3.248568880e-10 palpha0 = 4.930380658e-32
+ alpha1 = 0.0
+ beta0 = 1.443635041e+01 lbeta0 = 1.334731420e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.468709523e-01 lkt1 = -4.277743590e-8
+ kt2 = -3.564771813e-02 lkt2 = -2.847900921e-9
+ at = 6.717907755e+04 lat = -3.558108488e-2
+ ute = -1.241165273e+00 lute = 2.400093052e-7
+ ua1 = 1.881894468e-09 lua1 = 3.248571119e-16
+ ub1 = -1.042850307e-18 lub1 = -1.682422020e-24
+ uc1 = 1.351529876e-10 luc1 = -2.852147239e-16
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.67 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.293740921e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 9.044136365e-9
+ k1 = 4.583691775e-01 lk1 = -8.677927811e-10
+ k2 = -2.323755968e-02 lk2 = -9.089647275e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.295621900e+03 lvsat = 7.983307901e-2
+ ua = -7.179815791e-10 lua = -7.729276606e-16
+ ub = 2.353937299e-18 lub = 2.475523540e-25
+ uc = 5.823028540e-11 luc = -1.336786569e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.615025215e-02 lu0 = -9.319789778e-9
+ a0 = 2.215635936e+00 la0 = -7.186153452e-7
+ keta = -2.482972840e-01 lketa = 1.325215998e-07 wketa = -1.058791184e-22
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.193117478e+00 lags = 5.105707038e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.188839056e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.643919741e-9
+ nfactor = {7.336237045e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.168929469e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.487975000e-05 lcit = -9.642142013e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 5.649201940e-04 leta0 = -1.282790573e-10
+ etab = -5.274144355e-04 letab = 5.416955383e-11
+ dsub = 2.358547406e-01 ldsub = 3.287750393e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.565962295e-01 lpclm = -4.360176618e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 8.873827250e-03 lpdiblc2 = 5.679221645e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.999502351e-04 lalpha0 = -1.492145659e-10
+ alpha1 = 0.0
+ beta0 = 2.159946903e+01 lbeta0 = -8.066500302e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.675342905e-01 lkt1 = -1.947712687e-9
+ kt2 = -5.111828125e-02 lkt2 = 2.772115829e-8
+ at = 2.049761305e+04 lat = 5.665915489e-2
+ ute = -1.145855460e+00 lute = 5.168188119e-8
+ ua1 = 2.095780665e-09 lua1 = -9.777132001e-17
+ ub1 = -2.058942765e-18 lub1 = 3.253258715e-25
+ uc1 = 3.059635605e-11 luc1 = -7.861604784e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.68 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.468927403e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -8.053188390e-9
+ k1 = 4.428112210e-01 lk1 = 1.431599487e-8
+ k2 = -2.312855893e-02 lk2 = -9.196026549e-9
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.116988700e+02 lvsat = 8.128131369e-2
+ ua = -1.189585556e-09 lua = -3.126657592e-16
+ ub = 2.563393283e-18 lub = 4.313378596e-26
+ uc = 3.289414631e-11 luc = 1.135893926e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.043856181e-02 lu0 = -3.745465588e-9
+ a0 = 1.956396665e+00 la0 = -4.656107786e-7
+ keta = -2.196082690e-01 lketa = 1.045225556e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.134391582e+00 lags = -1.384015758e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.078412353e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -7.133174371e-9
+ nfactor = {1.560380996e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.620556907e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.733691026e-03 leta0 = 2.115050563e-09 weta0 = -4.135903063e-25 peta0 = 1.972152263e-31
+ etab = -8.021336290e-04 letab = 3.222817507e-10
+ dsub = 1.660149467e-01 ldsub = 3.969351861e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.044219330e-01 lpclm = 1.049127385e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.168699006e-02 lpdiblc2 = -6.825784599e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.221009338e-05 lalpha0 = 8.712180668e-11 palpha0 = -1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.743034605e+01 lbeta0 = 3.262205538e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.684353150e-01 lkt1 = -1.068357826e-9
+ kt2 = -1.026029230e-02 lkt2 = -1.215419603e-8
+ at = 7.584674830e+04 lat = 2.641166347e-3
+ ute = -1.058346030e+00 lute = -3.372294702e-8
+ ua1 = 2.504580930e-09 lua1 = -4.967399386e-16
+ ub1 = -2.138248650e-18 lub1 = 4.027244500e-25
+ uc1 = -8.636812690e-11 luc1 = 3.553543930e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.69 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955958815e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.123344844e-08 wvth0 = -2.117582368e-22
+ k1 = 3.575470440e-01 lk1 = 5.489747991e-8
+ k2 = -1.180429035e-02 lk2 = -1.458581218e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.920040959e+05 lvsat = -9.716707688e-3
+ ua = -1.540010971e-09 lua = -1.458807828e-16
+ ub = 2.620208842e-18 lub = 1.609242065e-26
+ uc = 7.025556412e-11 luc = -6.423227544e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.679655316e-02 lu0 = -2.012051571e-9
+ a0 = 4.931589960e-01 la0 = 2.308171899e-7
+ keta = 2.449876974e-02 lketa = -1.166018946e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.311916620e-01 lags = -9.742775603e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.329546542e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.819557388e-9
+ nfactor = {2.088047121e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.109129981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.810000000e-07 lcit = 2.150818050e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.566597539e-03 leta0 = 6.832822021e-11
+ etab = 7.541036029e-03 letab = -3.648649848e-09 wetab = 1.344168495e-24 petab = -7.642090019e-31
+ dsub = 1.588048920e+00 ldsub = -2.798818835e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.134240660e-01 lpclm = 1.006281733e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.854256280e-03 lpdiblc2 = 2.137655044e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.011350105e-03 lalpha0 = 5.483839952e-10 walpha0 = -2.067951531e-25 palpha0 = -2.465190329e-32
+ alpha1 = 0.0
+ beta0 = 1.918019144e+01 lbeta0 = 2.429366624e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701829100e-01 lkt1 = -2.365899855e-10
+ kt2 = -4.601988180e-02 lkt2 = 4.865580593e-9
+ at = 1.069337728e+05 lat = -1.215470296e-2
+ ute = -1.227804580e+00 lute = 4.693084985e-8
+ ua1 = 1.752556260e-09 lua1 = -1.388137969e-16
+ ub1 = -1.683418286e-18 lub1 = 1.862479382e-25 wub1 = 7.346839693e-40
+ uc1 = -2.881638008e-11 luc1 = 8.143685399e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.70 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.221476949e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.982783066e-8
+ k1 = 3.113341429e-01 lk1 = 6.533928492e-8
+ k2 = 2.363068596e-03 lk2 = -1.778692694e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.237662533e+05 lvsat = 5.701632855e-3
+ ua = -2.013580132e-09 lua = -3.887783096e-17
+ ub = 3.201343101e-18 lub = -1.152148652e-25
+ uc = 6.627162171e-11 luc = -5.523055757e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.577720036e-02 lu0 = -1.781728806e-9
+ a0 = 4.889235214e+00 la0 = -7.624762317e-7
+ keta = 1.417358112e-01 lketa = -3.814989897e-08 pketa = -6.310887242e-30
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.438389643e+00 lags = 5.509541398e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.642915643e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.190013221e-8
+ nfactor = {1.168008132e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 3.187958077e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 2.113928571e-05 lcit = -2.516921607e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.564206905e-01 leta0 = 3.599150595e-08 weta0 = 2.316105715e-23 peta0 = 5.522026337e-30
+ etab = 1.674259653e-02 letab = -5.727742443e-9
+ dsub = 3.726607961e-01 ldsub = -5.264936889e-9
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.261245636e+00 lpclm = -1.587221104e-7
+ pdiblc1 = -9.689928571e-01 lpdiblc1 = 3.070644361e-7
+ pdiblc2 = 7.663234286e-03 lpdiblc2 = 1.051066463e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.517701205e-03 lalpha0 = -4.749551482e-10
+ alpha1 = 0.0
+ beta0 = 3.347280247e+01 lbeta0 = -8.000488374e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.978221071e-01 lkt1 = -1.658651339e-8
+ kt2 = -3.256866571e-02 lkt2 = 1.826278318e-9
+ at = 6.586697143e+03 lat = 1.051871878e-2
+ ute = 6.271775714e-01 lute = -3.722023673e-7
+ ua1 = 4.205380043e-09 lua1 = -6.930293307e-16
+ ub1 = -3.760022786e-18 lub1 = 6.554567249e-25
+ uc1 = -4.836768571e-13 luc1 = 1.741911106e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.71 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 8.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.814329152e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -2.228836078e-08 wvth0 = 2.772986034e-08 pvth0 = -4.324471720e-15
+ k1 = 7.815716500e-01 lk1 = -7.994254317e-9
+ k2 = -1.596444210e-01 lk2 = 7.478141068e-09 wk2 = -8.910320961e-09 pk2 = 1.389564554e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.309759906e+05 lvsat = 4.577274319e-03 wvsat = 3.201821370e-02 pvsat = -4.993240427e-9
+ ua = -1.956579171e-09 lua = -4.776713090e-17 wua = -4.479281860e-17 pua = 6.985440061e-24
+ ub = 1.821001660e-18 lub = 1.000493826e-25 wub = 4.653091964e-25 pub = -7.256496917e-32
+ uc = 1.399819473e-10 luc = -1.701818103e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.072466544e-02 lu0 = -9.937859854e-10 wu0 = -6.069250387e-10 pu0 = 9.464995979e-17
+ a0 = 0.0
+ keta = 4.702508516e-01 lketa = -8.938181952e-08 wketa = -4.353714517e-07 pketa = 6.789617789e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.706276667e-01 lags = 9.729289038e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.105877863e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 3.525028035e-09 wvoff = 1.809103481e-12 pvoff = -2.821296878e-19
+ nfactor = {2.735001818e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 7.442314238e-08 wnfactor = -1.822097902e-06 pnfactor = 2.841561677e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.599166667e-05 lcit = 3.273650417e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.641077990e-01 leta0 = -2.958991198e-8
+ etab = -9.518338731e-02 letab = 1.172711474e-8
+ dsub = 6.699876640e-01 ldsub = -5.163306194e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -3.219917613e-01 lpclm = 8.818376168e-08 wpclm = 1.593178227e-07 ppclm = -2.484561444e-14
+ pdiblc1 = 1.0
+ pdiblc2 = -1.253275097e-02 lpdiblc2 = 4.200630363e-09 wpdiblc2 = 6.837633048e-09 ppdiblc2 = -1.066328874e-15
+ pdiblcb = 0.0
+ drout = -2.669909122e+01 ldrout = 4.708706146e-06 wdrout = 2.379262868e-05 pdrout = -3.710460443e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.391024405e-03 lalpha0 = -2.992499013e-10 walpha0 = 2.469620779e-11 palpha0 = -3.851373604e-18
+ alpha1 = 0.0
+ beta0 = 5.365279630e+01 lbeta0 = -3.947118875e-06 wbeta0 = 5.670469512e-06 pbeta0 = -8.843097205e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.219432500e-01 lkt1 = 1.836517884e-08 wkt1 = 1.361690792e-07 pkt1 = -2.123556790e-14
+ kt2 = -2.659712167e-02 lkt2 = 8.950160239e-10
+ at = 1.156654978e+05 lat = -6.492120182e-03 wat = -4.413823439e-02 pat = 6.883357653e-9
+ ute = -1.908540833e+00 lute = 2.324291796e-8
+ ua1 = -2.858552167e-10 lua1 = 7.378808039e-18
+ ub1 = 8.407201000e-19 lub1 = -6.202912810e-26
+ uc1 = -2.428191833e-11 luc1 = 5.453246864e-18
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.72 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.73 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {0.4229525+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = -0.057410608
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 200550.0
+ ua = -9.7927443e-10
+ ub = 2.30409e-18
+ uc = 2.2350587e-11
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 0.0312064
+ a0 = 1.9208155
+ keta = 0.0
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 0.537176
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6893098+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 0.08
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.2
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -0.25763
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.74 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.120860594e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.320442463e-8
+ k1 = 6.076841567e-01 lk1 = -2.959067260e-7
+ k2 = -8.662790178e-02 lk2 = 1.161664992e-07 wk2 = 5.293955920e-23
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.565038297e+05 lvsat = -6.200646292e-01 pvsat = 4.235164736e-22
+ ua = -8.509614041e-10 lua = -5.101661753e-16
+ ub = 2.131065938e-18 lub = 6.879350183e-25
+ uc = -6.413725184e-12 luc = 1.143654670e-16
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.098189256e-02 lu0 = 8.926303521e-10
+ a0 = 1.988847952e+00 la0 = -2.704936295e-7
+ keta = 1.790507093e-01 lketa = -7.118966674e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -3.661631337e-01 lags = 3.591631228e-6
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.035102483e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -2.673365840e-8
+ nfactor = {2.049039036e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -1.430265455e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 1.585440125e-01 leta0 = -3.122870665e-7
+ etab = -1.386642625e-01 letab = 2.730056745e-7
+ dsub = 7.158598930e-01 ldsub = -6.196911417e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.658852233e-01 lpclm = 1.356386466e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.440451272e-03 lpdiblc2 = 1.641530091e-8
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -3.997053919e-05 lalpha0 = 3.248568880e-10
+ alpha1 = 0.0
+ beta0 = 1.443635041e+01 lbeta0 = 1.334731420e-5
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.468709523e-01 lkt1 = -4.277743590e-8
+ kt2 = -3.564771813e-02 lkt2 = -2.847900921e-9
+ at = 6.717907755e+04 lat = -3.558108488e-2
+ ute = -1.241165272e+00 lute = 2.400093052e-7
+ ua1 = 1.881894467e-09 lua1 = 3.248571119e-16
+ ub1 = -1.042850307e-18 lub1 = -1.682422020e-24
+ uc1 = 1.351529876e-10 luc1 = -2.852147239e-16 puc1 = -9.403954807e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.75 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.135985294e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 2.378108594e-07 wvth0 = 6.807603084e-08 pvth0 = -1.345148331e-13
+ k1 = 5.783088781e-01 lk1 = -2.378626441e-07 wk1 = -7.052454393e-08 pk1 = 1.393529726e-13
+ k2 = -7.995537539e-02 lk2 = 1.029819207e-07 wk2 = 3.335007564e-08 pk2 = -6.589808197e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.314856358e+04 lvsat = -8.902911125e-04 wvsat = -2.402152971e-02 pvsat = 4.746534163e-8
+ ua = 1.037530780e-09 lua = -4.241732306e-15 wua = -1.032241267e-15 pua = 2.039657132e-21
+ ub = 2.144245332e-18 lub = 6.618931950e-25 wub = 1.232988762e-25 pub = -2.436324145e-31
+ uc = -4.622147905e-11 luc = 1.930235983e-16 wuc = 6.141763749e-17 puc = -1.213581808e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 5.747911668e-02 lu0 = -5.146455965e-08 wu0 = -1.254137234e-08 pu0 = 2.478112468e-14
+ a0 = 2.650291794e+00 la0 = -1.577473589e-06 wa0 = -2.555776448e-07 pa0 = 5.050086473e-13
+ keta = -3.427477731e-01 lketa = 3.191510438e-07 wketa = 5.553688759e-08 pketa = -1.097381130e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 1.422250368e+00 lags = 5.781556913e-08 wags = -1.347301395e-07 pags = 2.662200192e-13
+ b0 = 4.353092896e-07 lb0 = -8.601493909e-13 wb0 = -2.559618623e-13 pb0 = 5.057678418e-19
+ b1 = 1.199991034e-08 lb1 = -2.371122283e-14 wb1 = -7.055947279e-15 pb1 = 1.394219903e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.999238293e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.637747570e-07 wvoff = 4.765147514e-08 pvoff = -9.415693231e-14
+ nfactor = {-1.998211804e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 6.566899841e-06 wnfactor = 1.606319279e-06 pnfactor = -3.174006579e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.188103333e-05 lcit = -6.299532782e-11 wcit = -1.587675460e-11 pcit = 3.137167325e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.429567401e-03 leta0 = 3.812728706e-09 weta0 = 1.172758706e-09 peta0 = -2.317312565e-15
+ etab = 2.021020688e-03 letab = -4.981410829e-09 wetab = -1.498479853e-09 petab = 2.960921265e-15
+ dsub = -1.452976545e+00 ldsub = 3.665821218e-06 wdsub = 9.930327960e-07 pdsub = -1.962183153e-12
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 4.313485352e-01 lpclm = -3.889035847e-07 wpclm = -1.027543558e-07 ppclm = 2.030374693e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -8.450196137e-03 lpdiblc2 = 3.991062566e-08 wpdiblc2 = 1.018652575e-08 ppdiblc2 = -2.012806556e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.232495306e-04 lalpha0 = -5.904428088e-10 walpha0 = -1.312999858e-10 palpha0 = 2.594422069e-16
+ alpha1 = 0.0
+ beta0 = 2.769130957e+01 lbeta0 = -1.284382234e-05 wbeta0 = -3.582002236e-06 pbeta0 = 7.077857317e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -1.919846997e-01 lkt1 = -1.512299266e-07 wkt1 = -4.442315937e-08 pkt1 = 8.777794176e-14
+ kt2 = -9.992580100e-02 lkt2 = 1.241623769e-07 wkt2 = 2.869882161e-08 pkt2 = -5.670743657e-14
+ at = 5.553987856e+04 lat = -1.258260964e-02 wat = -2.060485212e-02 pat = 4.071415755e-8
+ ute = -9.487460917e-01 lute = -3.377963752e-07 wute = -1.159003086e-07 pute = 2.290132147e-13
+ ua1 = 2.702769514e-09 lua1 = -1.297150937e-15 wua1 = -3.569094434e-16 pua1 = 7.052352147e-22
+ ub1 = -2.981846629e-18 lub1 = 2.148937762e-24 wub1 = 5.426674722e-25 pub1 = -1.072283792e-30
+ uc1 = 5.046686881e-10 luc1 = -1.015359272e-15 wuc1 = -2.787545312e-16 puc1 = 5.508050160e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.76 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {6.784438656e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.182599465e-07 wvth0 = -1.361520617e-07 pvth0 = 6.480157376e-14
+ k1 = 2.029318199e-01 lk1 = 1.284865958e-07 wk1 = 1.410490879e-07 pk1 = -6.713231337e-14
+ k2 = 9.030707250e-02 lk2 = -6.318571533e-08 wk2 = -6.670015129e-08 pk2 = 3.174593700e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -8.089418450e+04 lvsat = 1.201692289e-01 wvsat = 4.804305942e-02 pvsat = -2.286609413e-8
+ ua = -4.700610274e-09 lua = 1.358406455e-15 wua = 2.064482534e-15 pua = -9.825904622e-22
+ ub = 2.982777216e-18 lub = -1.564719968e-25 wub = -2.465977524e-25 pub = 1.173682003e-31
+ uc = 2.417976752e-10 luc = -8.806869531e-17 wuc = -1.228352750e-16 puc = 5.846344913e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -1.221916726e-02 lu0 = 1.655748056e-08 wu0 = 2.508274469e-08 pu0 = -1.193813233e-14
+ a0 = 1.087084948e+00 la0 = -5.186186682e-08 wa0 = 5.111552897e-07 pa0 = -2.432843601e-13
+ keta = -3.070729080e-02 lketa = 1.461513506e-08 wketa = -1.110737752e-07 pketa = 5.286556330e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 2.676125801e+00 lags = -1.165904160e-06 wags = 2.694602791e-07 pags = -1.282496198e-13
+ b0 = -8.706185793e-07 lb0 = 4.143709128e-13 wb0 = 5.119237246e-13 pb0 = -2.436500967e-19
+ b1 = -2.399982068e-08 lb1 = 1.142271465e-14 wb1 = 1.411189456e-14 pb1 = -6.716556215e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {5.423861216e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -8.427507775e-08 wvoff = -9.530295029e-08 pvoff = 4.535943919e-14
+ nfactor = {7.024052012e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -2.238378530e-06 wnfactor = -3.212638558e-06 pnfactor = 1.529055322e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -4.900256667e-05 lcit = 2.570252161e-11 wcit = 3.175350920e-11 pcit = -1.511308270e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.255284165e-03 leta0 = 2.164978206e-10 weta0 = -2.345517412e-09 peta0 = 1.116349012e-15
+ etab = -5.899003876e-03 letab = 2.748137145e-09 wetab = 2.996959705e-09 petab = -1.426402972e-15
+ dsub = 3.543677518e+00 ldsub = -1.210663315e-06 wdsub = -1.986065592e-06 pdsub = 9.452679186e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -2.450826785e-01 lpclm = 2.712594583e-07 wpclm = 2.055087115e-07 ppclm = -9.781187126e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 5.633503683e-02 lpdiblc2 = -2.331652246e-08 wpdiblc2 = -2.037305150e-08 ppdiblc2 = 9.696553863e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.888086844e-04 lalpha0 = 2.996804061e-10 walpha0 = 2.625999715e-10 palpha0 = -1.249844564e-16
+ alpha1 = 0.0
+ beta0 = 5.246664980e+00 lbeta0 = 9.061028545e-06 wbeta0 = 7.164004471e-06 pbeta0 = -3.409707928e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -4.195344965e-01 lkt1 = 7.084729763e-08 wkt1 = 8.884631874e-08 pkt1 = -4.228640541e-14
+ kt2 = 8.735474721e-02 lkt2 = -5.861407408e-08 wkt2 = -5.739764323e-08 pkt2 = 2.731840830e-14
+ at = 5.762217280e+03 lat = 3.599789889e-02 wat = 4.120970424e-02 pat = -1.961375873e-8
+ ute = -1.452564767e+00 lute = 1.539054607e-07 wute = 2.318006172e-07 pute = -1.103255037e-13
+ ua1 = 1.290603231e-09 lua1 = 8.105274705e-17 wua1 = 7.138188868e-16 pua1 = -3.397420992e-22
+ ub1 = -2.924409213e-19 lub1 = -4.757877385e-25 wub1 = -1.085334944e-24 pub1 = 5.165651668e-31
+ uc1 = -1.034512791e-09 luc1 = 4.868048921e-16 wuc1 = 5.575090624e-16 puc1 = -2.653464383e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.77 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955958815e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.123344844e-8
+ k1 = 3.575470440e-01 lk1 = 5.489747991e-8
+ k2 = -1.180429035e-02 lk2 = -1.458581218e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.920040959e+05 lvsat = -9.716707688e-3
+ ua = -1.540010971e-09 lua = -1.458807828e-16
+ ub = 2.620208842e-18 lub = 1.609242065e-26
+ uc = 7.025556412e-11 luc = -6.423227544e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.679655316e-02 lu0 = -2.012051571e-9
+ a0 = 4.931589960e-01 la0 = 2.308171899e-7
+ keta = 2.449876974e-02 lketa = -1.166018946e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.311916620e-01 lags = -9.742775603e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.329546542e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.819557388e-9
+ nfactor = {2.088047121e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.109129981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.810000000e-07 lcit = 2.150818050e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.566597539e-03 leta0 = 6.832822021e-11
+ etab = 7.541036029e-03 letab = -3.648649848e-09 wetab = 1.344168495e-24 petab = -6.162975822e-31
+ dsub = 1.588048920e+00 ldsub = -2.798818835e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.134240660e-01 lpclm = 1.006281733e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.854256280e-03 lpdiblc2 = 2.137655044e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.011350105e-03 lalpha0 = 5.483839952e-10 walpha0 = -1.033975766e-25 palpha0 = -1.479114197e-31
+ alpha1 = 0.0
+ beta0 = 1.918019144e+01 lbeta0 = 2.429366624e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701829100e-01 lkt1 = -2.365899855e-10
+ kt2 = -4.601988180e-02 lkt2 = 4.865580593e-09 wkt2 = -2.646977960e-23
+ at = 1.069337728e+05 lat = -1.215470296e-2
+ ute = -1.227804580e+00 lute = 4.693084985e-08 wute = 8.470329473e-22
+ ua1 = 1.752556260e-09 lua1 = -1.388137969e-16
+ ub1 = -1.683418286e-18 lub1 = 1.862479382e-25
+ uc1 = -2.881638008e-11 luc1 = 8.143685399e-18 puc1 = -2.938735877e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.78 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {1.210981923e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -1.928749244e-07 wvth0 = -3.462345259e-07 pvth0 = 7.823169113e-14
+ k1 = -1.703003519e-01 lk1 = 1.741645990e-07 wk1 = 2.832010829e-07 pk1 = -6.398928469e-14
+ k2 = 1.528862373e-01 lk2 = -5.179763691e-08 wk2 = -8.850762321e-08 pk2 = 1.999829746e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.323461767e+05 lvsat = 3.762999156e-03 wvsat = -5.044994976e-03 pvsat = 1.139916615e-9
+ ua = 3.779380764e-09 lua = -1.347797345e-15 wua = -3.406261007e-15 pua = 7.696446744e-22
+ ub = 5.006338575e-18 lub = -5.230535926e-25 wub = -1.061337339e-24 pub = 2.398091717e-31
+ uc = -2.331315495e-10 luc = 6.212709077e-17 wuc = 1.760490646e-16 puc = -3.977828616e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 1.215349397e-01 lu0 = -2.341819002e-08 wu0 = -5.630555075e-08 pu0 = 1.272223919e-14
+ a0 = 4.889235214e+00 la0 = -7.624762317e-7
+ keta = 1.410149654e+00 lketa = -3.247480068e-07 wketa = -7.458273397e-07 pketa = 1.685196874e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.377985010e+00 lags = 5.373057129e-07 wags = -3.551792440e-08 pags = 8.025275018e-15
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-5.870528927e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.074230544e-07 wvoff = 2.485836611e-07 pvoff = -5.616747823e-14
+ nfactor = {-4.185855458e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.528501286e-06 wnfactor = 3.148071791e-06 pnfactor = -7.113068212e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 8.277666667e-05 lcit = -1.644388783e-11 wcit = -3.624278000e-11 pcit = 8.189056141e-18
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.772218519e-01 leta0 = 4.069152838e-08 weta0 = 1.223108292e-08 peta0 = -2.763613186e-15
+ etab = -1.239928766e-01 letab = 2.607143771e-08 wetab = 8.275245821e-08 petab = -1.869791793e-14
+ dsub = 1.161827230e-01 ldsub = 5.268628374e-08 wdsub = 1.508091070e-07 pdsub = -3.407531773e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 2.096062323e+00 lpclm = -3.473489410e-07 wpclm = -4.908722123e-07 ppclm = 1.109125764e-13
+ pdiblc1 = -1.281569748e+01 lpdiblc1 = 2.983827345e-06 wpdiblc1 = 6.965862316e-06 ppdiblc1 = -1.573936590e-12
+ pdiblc2 = -1.773136667e-02 lpdiblc2 = 6.788976548e-09 wpdiblc2 = 1.493202536e-08 ppdiblc2 = -3.373891130e-15
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.916425163e-03 lalpha0 = -5.650468265e-10 walpha0 = -2.344496873e-10 palpha0 = 5.297390684e-17
+ alpha1 = 0.0
+ beta0 = 3.660108447e+01 lbeta0 = -1.506884154e-06 wbeta0 = -1.839429813e-06 pbeta0 = 4.156191663e-13
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = 2.351188567e-01 lkt1 = -1.144095242e-07 wkt1 = -2.545692867e-07 pkt1 = 5.751993033e-14
+ kt2 = -1.447117166e-01 lkt2 = 2.716500067e-08 wkt2 = 6.594011393e-08 pkt2 = -1.489916874e-14
+ at = -4.649541533e+04 lat = 2.251262209e-02 wat = 3.121228214e-02 pat = -7.052415149e-9
+ ute = 8.466066476e-01 lute = -4.217823670e-07 wute = -1.290242968e-07 pute = 2.915303986e-14
+ ua1 = 6.131918022e-09 lua1 = -1.128330587e-15 wua1 = -1.132804332e-15 pua1 = 2.559571387e-22
+ ub1 = -6.905008511e-18 lub1 = 1.366066250e-24 wub1 = 1.849251607e-24 pub1 = -4.178384005e-31
+ uc1 = -2.032164193e-10 luc1 = 4.754937426e-17 wuc1 = 1.192068526e-16 puc1 = -2.693478833e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.79 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 6.4e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.024292173e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 1.557160707e-07 wvth0 = 8.542962120e-07 pvth0 = -1.089910774e-13
+ k1 = 1.905385471e+00 lk1 = -1.495386051e-07 wk1 = -6.608025268e-07 pk1 = 8.322807825e-14
+ k2 = -5.045140241e-01 lk2 = 5.072393386e-08 wk2 = 1.938730057e-07 pk2 = -2.403896161e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.035329431e+05 lvsat = -7.338577058e-03 wvsat = -1.064527435e-02 pvsat = 2.013280183e-9
+ ua = -1.439916192e-08 lua = 1.487146386e-15 wua = 7.271445838e-15 pua = -8.955437080e-22
+ ub = 1.500370403e-18 lub = 2.370214389e-26 wub = 6.538403753e-25 pub = -2.767279281e-32
+ uc = 1.387267795e-09 luc = -1.905741870e-16 wuc = -7.334040783e-16 puc = 1.020509315e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = -2.018930753e-01 lu0 = 2.702040893e-08 wu0 = 1.302923065e-07 pu0 = -1.637769665e-14
+ a0 = 0.0
+ keta = -3.228694010e+00 lketa = 3.986796627e-07 wketa = 1.739608127e-06 pketa = -2.190839736e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.296835222e-01 lags = 1.150448054e-07 wags = 8.287515693e-08 pags = -1.043812602e-14
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {8.758816209e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.207215830e-07 wvoff = -5.800422023e-07 pvoff = 7.305672517e-14
+ nfactor = {8.258296662e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -4.121642373e-07 wnfactor = -5.069795270e-06 pnfactor = 5.702695470e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -1.598122222e-04 lcit = 2.138784939e-11 wcit = 8.456648667e-11 pcit = -1.065114900e-17
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.126438423e-01 leta0 = -3.570302664e-08 weta0 = -2.853919348e-08 peta0 = 3.594511419e-15
+ etab = 2.331993834e-01 letab = -2.963269523e-08 wetab = -1.930890692e-07 petab = 2.431956826e-14
+ dsub = 1.268436501e+00 ldsub = -1.270076930e-07 wdsub = -3.518879163e-07 pdsub = 4.432028306e-14
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -7.763128533e-01 lpclm = 1.005979678e-07 wpclm = 4.264586248e-07 ppclm = -3.214516767e-14
+ pdiblc1 = 2.864231078e+01 lpdiblc1 = -3.481549042e-06 wpdiblc1 = -1.625367874e-05 ppdiblc1 = 2.047150837e-12
+ pdiblc2 = -8.867764700e-02 lpdiblc2 = 1.785304897e-08 wpdiblc2 = 5.161083192e-08 ppdiblc2 = -9.093951013e-15
+ pdiblcb = 0.0
+ drout = 7.059169160e+01 ldrout = -1.046379144e-05 wdrout = -3.341435162e-05 pdrout = 5.210968135e-12
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 1.452065253e-03 lalpha0 = -1.807298987e-10 walpha0 = 5.768041890e-10 palpha0 = -7.354113517e-17
+ alpha1 = 0.0
+ beta0 = 3.153511828e+01 lbeta0 = -7.168467270e-07 wbeta0 = 1.867566419e-05 pbeta0 = -2.783709743e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -8.753278767e-01 lkt1 = 5.876464390e-08 wkt1 = 4.027592397e-07 pkt1 = -4.499045336e-14
+ kt2 = 2.350699971e-01 lkt2 = -3.206195759e-08 wkt2 = -1.538602658e-07 pkt2 = 1.937870048e-14
+ at = 2.320835299e+05 lat = -2.093176441e-02 wat = -1.125920373e-01 pat = 1.537386846e-8
+ ute = -2.420542011e+00 lute = 8.772946630e-08 wute = 3.010566925e-07 pute = -3.791809042e-14
+ ua1 = -7.315356049e-09 lua1 = 9.687718043e-16 wua1 = 4.133346489e-15 pua1 = -5.652990818e-22
+ ub1 = 8.179020127e-18 lub1 = -9.862880165e-25 wub1 = -4.314920416e-24 pub1 = 5.434642264e-31
+ uc1 = 4.487611474e-10 luc1 = -5.412652726e-17 wuc1 = -2.781493226e-16 puc1 = 3.503290718e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.80 nmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.392302723e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = -8.106330609e-9
+ k1 = 6.849043077e-01 wk1 = -7.551886523e-8
+ k2 = -9.805085218e-02 wk2 = 2.023884160e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.087896308e+05 wvsat = -1.535033361e-1
+ ua = -3.972615672e-10 wua = -2.898424057e-16
+ ub = 1.554870308e-18 wub = 3.731114068e-25
+ uc = 1.431003328e-11 wuc = 4.004195754e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.306338462e-02 wu0 = -9.247783385e-10
+ a0 = 2.942767069e+00 wa0 = -5.089318815e-7
+ keta = 3.680000000e-01 wketa = -1.832640000e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.920676554e+00 wags = 1.722010572e-6
+ b0 = -2.281854769e-07 wb0 = 1.136363675e-13
+ b1 = -6.290252308e-09 wb1 = 3.132545649e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-5.383729738e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = -2.808560272e-8
+ nfactor = {2.436130472e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -3.719166947e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.062799503e-01 weta0 = -1.126874152e-7
+ etab = -2.681538462e-01 wetab = 9.868061538e-8
+ dsub = 1.409230769e+00 wdsub = -4.229169231e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 7.465353846e-02 wpclm = 6.242253785e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -3.515909231e-03 wpdiblc2 = 5.520334597e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.038681500e-05 walpha0 = 6.579663250e-11
+ alpha1 = 0.0
+ beta0 = 6.165573585e+00 wbeta0 = 5.790639129e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.635463077e-01 wkt1 = 2.946321231e-9
+ kt2 = -4.941950769e-02 wkt2 = 6.501642831e-9
+ at = -1.766858462e+04 wat = 3.779749514e-2
+ ute = -1.532947692e+00 wute = 1.753695508e-7
+ ua1 = 1.554836923e-09 wua1 = 2.035640123e-16
+ ub1 = -2.473538462e-19 wub1 = -6.068857846e-25
+ uc1 = 1.358517231e-10 wuc1 = -3.607199409e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.81 nmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.392302723e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = -8.106330609e-9
+ k1 = 6.849043077e-01 wk1 = -7.551886523e-8
+ k2 = -9.805085218e-02 wk2 = 2.023884160e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.087896308e+05 wvsat = -1.535033361e-1
+ ua = -3.972615672e-10 wua = -2.898424057e-16
+ ub = 1.554870308e-18 wub = 3.731114068e-25
+ uc = 1.431003328e-11 wuc = 4.004195754e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.306338462e-02 wu0 = -9.247783385e-10
+ a0 = 2.942767069e+00 wa0 = -5.089318815e-7
+ keta = 3.680000000e-01 wketa = -1.832640000e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.920676554e+00 wags = 1.722010572e-6
+ b0 = -2.281854769e-07 wb0 = 1.136363675e-13
+ b1 = -6.290252308e-09 wb1 = 3.132545649e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-5.383729738e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} wvoff = -2.808560272e-8
+ nfactor = {2.436130472e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -3.719166947e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.062799503e-01 weta0 = -1.126874152e-7
+ etab = -2.681538462e-01 wetab = 9.868061538e-8
+ dsub = 1.409230769e+00 wdsub = -4.229169231e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 7.465353846e-02 wpclm = 6.242253785e-8
+ pdiblc1 = 0.39
+ pdiblc2 = -3.515909231e-03 wpdiblc2 = 5.520334597e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -9.038681500e-05 walpha0 = 6.579663250e-11
+ alpha1 = 0.0
+ beta0 = 6.165573585e+00 wbeta0 = 5.790639129e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.635463077e-01 wkt1 = 2.946321231e-9
+ kt2 = -4.941950769e-02 wkt2 = 6.501642831e-9
+ at = -1.766858462e+04 wat = 3.779749514e-2
+ ute = -1.532947692e+00 wute = 1.753695508e-7
+ ua1 = 1.554836923e-09 wua1 = 2.035640123e-16
+ ub1 = -2.473538462e-19 wub1 = -6.068857846e-25
+ uc1 = 1.358517231e-10 wuc1 = -3.607199409e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.82 nmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {3.976034459e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.655061805e-07 wvth0 = 7.212341514e-09 pvth0 = -6.090627443e-14
+ k1 = 9.700060774e-01 lk1 = -1.133550381e-06 wk1 = -1.804363165e-07 pk1 = 4.171465403e-13
+ k2 = -2.099755622e-01 lk2 = 4.450070508e-07 wk2 = 6.142713489e-08 pk2 = -1.637625947e-13
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.106212763e+06 lvsat = -2.375324503e+00 wvsat = -3.733550488e-01 pvsat = 8.741194170e-7
+ ua = 9.427602426e-11 lua = -1.954328887e-15 wua = -4.707282393e-16 pua = 7.191930304e-22
+ ub = 8.920550558e-19 lub = 2.635320301e-24 wub = 6.170274195e-25 pub = -9.697978707e-31
+ uc = -9.587940878e-11 luc = 4.381077121e-16 wuc = 4.455391043e-17 puc = -1.612236381e-22
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.220334843e-02 lu0 = 3.419460887e-09 wu0 = -6.082850208e-10 pu0 = -1.258361607e-15
+ a0 = 3.203383695e+00 la0 = -1.036198673e-06 wa0 = -6.048387997e-07 pa0 = 3.813211116e-13
+ keta = 1.053901948e+00 lketa = -2.727111849e-06 wketa = -4.356759168e-07 pketa = 1.003577160e-12
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -6.381160312e+00 lags = 1.375871040e-05 wags = 2.995468595e-06 pags = -5.063205427e-12
+ b0 = -2.281854769e-07 wb0 = 1.136363675e-13
+ b1 = -6.290252308e-09 wb1 = 3.132545649e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.807981150e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.024104760e-07 wvoff = -3.756435753e-08 pvoff = 3.768705518e-14
+ nfactor = {3.814170160e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -5.479016896e-06 wnfactor = -8.790352997e-07 pnfactor = 2.016278218e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 6.071639366e-01 leta0 = -1.196299686e-06 weta0 = -2.234127222e-07 peta0 = 4.402382843e-13
+ etab = -5.311907902e-01 letab = 1.045821738e-06 wetab = 1.954782108e-07 petab = -3.848623995e-13
+ dsub = 2.006294052e+00 ldsub = -2.373893758e-06 wdsub = -6.426362111e-07 pdsub = 8.735929030e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.603229863e-02 lpclm = 5.196003540e-07 wpclm = 1.105149259e-07 ppclm = -1.912129303e-13
+ pdiblc1 = 0.39
+ pdiblc2 = -1.933180974e-02 lpdiblc2 = 6.288322963e-08 wpdiblc2 = 1.134058598e-08 ppdiblc2 = -2.314102850e-14
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -4.033816392e-04 lalpha0 = 1.244451771e-09 walpha0 = 1.809787278e-10 palpha0 = -4.579582518e-16
+ alpha1 = 0.0
+ beta0 = -6.694366949e+00 lbeta0 = 5.113048057e-05 wbeta0 = 1.052309725e-05 pbeta0 = -1.881601685e-11
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.223308786e-01 lkt1 = -1.638704852e-07 wkt1 = -1.222095667e-08 pkt1 = 6.030433856e-14
+ kt2 = -4.667559712e-02 lkt2 = -1.090965122e-08 wkt2 = 5.491883742e-09 pkt2 = 4.014751649e-15
+ at = 1.661326631e+04 lat = -1.363029252e-01 wat = 2.518177400e-02 pat = 5.015947646e-8
+ ute = -1.764193121e+00 lute = 9.194202614e-07 wute = 2.604678685e-07 pute = -3.383466562e-13
+ ua1 = 1.241841883e-09 lua1 = 1.244452629e-15 wua1 = 3.187461870e-16 pua1 = -4.579585674e-22
+ ub1 = 1.373634976e-18 lub1 = -6.444970507e-24 wub1 = -1.203409671e-24 pub1 = 2.371749147e-30
+ uc1 = 4.106519063e-10 luc1 = -1.092591789e-15 wuc1 = -1.371984615e-16 puc1 = 4.020737782e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.83 nmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.439822223e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.237309628e-07 wvth0 = -4.665504821e-08 pvth0 = 4.553299431e-14
+ k1 = 3.149796719e-01 lk1 = 1.607490447e-07 wk1 = 6.061340075e-08 pk1 = -5.915564846e-14
+ k2 = 7.212438997e-02 lk2 = -1.124083497e-07 wk2 = -4.238564751e-08 pk2 = 4.136627269e-14
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.789599465e+05 lvsat = 3.617075127e-01 wvsat = 1.363885083e-01 pvsat = -1.331083647e-7
+ ua = -6.116636638e-10 lua = -5.594273603e-16 wua = -2.109424341e-16 pua = 2.058692686e-22
+ ub = 1.890995166e-18 lub = 6.614645894e-25 wub = 2.494174588e-25 pub = -2.434189689e-31
+ uc = 2.240696379e-10 luc = -1.940956067e-16 wuc = -7.318733875e-17 puc = 7.142718326e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.723600433e-02 lu0 = -6.524815545e-09 wu0 = -2.460302393e-09 pu0 = 2.401132121e-15
+ a0 = 3.771240529e+00 la0 = -2.158255384e-06 wa0 = -8.138101147e-07 pa0 = 7.942379814e-13
+ keta = -5.177807955e-01 lketa = 3.784546674e-07 wketa = 1.427033327e-07 pketa = -1.392713176e-13
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -5.665465853e-01 lags = 2.269324405e-06 wags = 8.556907434e-07 pags = -8.351113810e-13
+ b0 = -5.295534467e-07 lb0 = 5.954880398e-13 wb0 = 2.245397804e-13 pb0 = -2.191395987e-19
+ b1 = -1.459788254e-08 lb1 = 1.641546196e-14 wb1 = 6.189753576e-15 pb1 = -6.040890002e-21
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-3.086818227e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -9.690079479e-08 wvoff = -3.653823708e-08 pvoff = 3.565949248e-14
+ nfactor = {6.663883198e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 7.408426302e-07 wnfactor = 2.793484174e-07 pnfactor = -2.726300879e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 3.363289817e-03 leta0 = -3.219797456e-09 weta0 = -1.214084189e-09 peta0 = 1.184885464e-15
+ etab = -3.784704231e-03 letab = 3.693682094e-09 wetab = 1.392771157e-09 petab = -1.359275011e-15
+ dsub = 1.336695973e+00 ldsub = -1.050801435e-06 wdsub = -3.962241182e-07 pdsub = 3.866949281e-13
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.704782675e-01 lpclm = 7.202680083e-08 wpclm = 2.715903756e-08 ppclm = -2.650586271e-14
+ pdiblc1 = 0.39
+ pdiblc2 = 1.347575443e-02 lpdiblc2 = -1.942876781e-09 wpdiblc2 = -7.325976285e-10 ppdiblc2 = 7.149786556e-16
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.611076608e-04 lalpha0 = -2.661408611e-10 walpha0 = -1.003533346e-10 palpha0 = 9.793983690e-17
+ alpha1 = 0.0
+ beta0 = 1.652845939e+01 lbeta0 = 5.243336867e-06 wbeta0 = 1.977097154e-06 pbeta0 = -1.929547967e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -3.537909218e-01 lkt1 = 9.588798716e-08 wkt1 = 3.615633923e-08 pkt1 = -3.528677928e-14
+ kt2 = -7.214993296e-02 lkt2 = 3.942636267e-08 wkt2 = 1.486643933e-08 pkt2 = -1.450890146e-14
+ at = -1.864726815e+05 lat = 2.649847534e-01 wat = 9.991740280e-02 pat = -9.751438926e-8
+ ute = -1.535543556e+00 lute = 4.676201531e-07 wute = 1.763248285e-07 pute = -1.720842163e-13
+ ua1 = 1.640967498e-09 lua1 = 4.558003704e-16 wua1 = 1.718679608e-16 pua1 = -1.677345363e-22
+ ub1 = -1.879847301e-18 lub1 = -1.625220121e-26 wub1 = -6.128193090e-27 pub1 = 5.980810047e-33
+ uc1 = -3.180843428e-10 luc1 = 3.473546029e-16 wuc1 = 1.309764782e-16 puc1 = -1.278264939e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.84 nmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.050461514e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.186369560e-8
+ k1 = 4.861629200e-01 lk1 = -6.317246274e-9
+ k2 = -4.362897425e-02 lk2 = 5.611461224e-10 wk2 = -1.323488980e-23
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.557782237e+04 lvsat = 7.425337721e-2
+ ua = -5.550630167e-10 lua = -6.146667619e-16
+ ub = 2.487601006e-18 lub = 7.920712019e-26
+ uc = -4.859503495e-12 luc = 2.932778889e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 3.814778995e-02 lu0 = -7.414672723e-9
+ a0 = 2.113501192e+00 la0 = -5.403846783e-7
+ keta = -2.537470000e-01 lketa = 1.207708847e-7
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 3.217210699e+00 lags = -1.423433517e-6
+ b0 = 1.573407071e-07 lb0 = -7.488630954e-14
+ b1 = 4.337316990e-09 lb1 = -2.064346021e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.371327740e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 6.808133470e-9
+ nfactor = {5.729705708e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 8.320136823e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.475950000e-05 lcit = -4.645034025e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -2.454590156e-03 leta0 = 2.458162504e-09 weta0 = -1.033975766e-25 peta0 = -1.109335648e-31
+ etab = 1.189875000e-04 letab = -1.161258506e-10
+ dsub = -4.444060000e-01 ldsub = 6.874650357e-07 pdsub = 5.048709793e-29
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.675854170e-01 lpclm = 7.485007828e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.542529486e-02 lpdiblc2 = -3.845530769e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.850049536e-05 lalpha0 = 4.870760197e-11
+ alpha1 = 0.0
+ beta0 = 1.963221613e+01 lbeta0 = 2.214225476e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.411282340e-01 lkt1 = -1.406516303e-8
+ kt2 = -2.790156450e-02 lkt2 = -3.757832526e-9
+ at = 8.851262740e+04 lat = -3.387158811e-3
+ ute = -9.871016800e-01 lute = -6.763169540e-8
+ ua1 = 2.723974490e-09 lua1 = -6.011603035e-16
+ ub1 = -2.471828360e-18 lub1 = 5.614917129e-25
+ uc1 = 8.498331840e-11 luc1 = -4.601928109e-17 wuc1 = 1.232595164e-32 puc1 = 5.877471754e-39
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.85 nmos
* DC IV MOS Parameters
+ lmin = 2.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {4.955958815e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -3.123344844e-8
+ k1 = 3.575470440e-01 lk1 = 5.489747991e-8
+ k2 = -1.180429035e-02 lk2 = -1.458581218e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.920040959e+05 lvsat = -9.716707688e-3
+ ua = -1.540010971e-09 lua = -1.458807828e-16
+ ub = 2.620208842e-18 lub = 1.609242065e-26
+ uc = 7.025556412e-11 luc = -6.423227544e-18
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 2.679655316e-02 lu0 = -2.012051571e-9
+ a0 = 4.931589960e-01 la0 = 2.308171899e-7
+ keta = 2.449876974e-02 lketa = -1.166018946e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.311916620e-01 lags = -9.742775603e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.329546542e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.819557388e-9
+ nfactor = {2.088047121e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.109129981e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 4.810000000e-07 lcit = 2.150818050e-12
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.566597539e-03 leta0 = 6.832822021e-11
+ etab = 7.541036029e-03 letab = -3.648649848e-09 wetab = 3.101927297e-25 petab = -2.465190329e-31
+ dsub = 1.588048920e+00 ldsub = -2.798818835e-7
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.134240660e-01 lpclm = 1.006281733e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.854256280e-03 lpdiblc2 = 2.137655044e-9
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = -1.011350105e-03 lalpha0 = 5.483839952e-10 walpha0 = -5.169878828e-26 palpha0 = 1.232595164e-32
+ alpha1 = 0.0
+ beta0 = 1.918019144e+01 lbeta0 = 2.429366624e-6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.701829100e-01 lkt1 = -2.365899855e-10
+ kt2 = -4.601988180e-02 lkt2 = 4.865580593e-9
+ at = 1.069337728e+05 lat = -1.215470296e-2
+ ute = -1.227804580e+00 lute = 4.693084985e-8
+ ua1 = 1.752556260e-09 lua1 = -1.388137969e-16
+ ub1 = -1.683418286e-18 lub1 = 1.862479382e-25
+ uc1 = -2.881638008e-11 luc1 = 8.143685399e-18 wuc1 = -6.162975822e-33
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.86 nmos
* DC IV MOS Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {5.157318706e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -3.578317517e-8
+ k1 = 3.983765214e-01 lk1 = 4.567205948e-8
+ k2 = -2.483991370e-02 lk2 = -1.164041308e-8
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.222156647e+05 lvsat = 6.051988343e-3
+ ua = -3.060500776e-09 lua = 1.976738885e-16
+ ub = 2.875139100e-18 lub = -4.150907114e-26
+ uc = 1.203806285e-10 luc = -1.774898585e-17
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 8.471584807e-03 lu0 = 2.128475028e-9
+ a0 = 4.889235214e+00 la0 = -7.624762317e-7
+ keta = -8.749560622e-02 lketa = 1.364493979e-8
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = -2.449306143e+00 lags = 5.534207230e-7
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.788891456e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -5.363046493e-9
+ nfactor = {2.135573841e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.001743357e-7
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = -1.526614445e-01 leta0 = 3.514210431e-08 weta0 = -9.926167351e-24
+ etab = 4.217671818e-02 letab = -1.147458223e-08 petab = 7.888609052e-31
+ dsub = 4.190122551e-01 ldsub = -1.573804905e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 1.110375150e+00 lpclm = -1.246329241e-7
+ pdiblc1 = 1.171977857e+00 lpdiblc1 = -1.766878968e-7
+ pdiblc2 = 1.225262000e-02 lpdiblc2 = 1.409476100e-11
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.445642658e-03 lalpha0 = -4.586735196e-10
+ alpha1 = 0.0
+ beta0 = 3.290745030e+01 lbeta0 = -6.723075151e-7
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -2.760644500e-01 lkt1 = 1.092343977e-9
+ kt2 = -1.230184929e-02 lkt2 = -2.753008854e-9
+ at = 1.617985000e+04 lat = 8.351145893e-3
+ ute = 5.875217143e-01 lute = -3.632421263e-7
+ ua1 = 3.857210529e-09 lua1 = -6.143604289e-16
+ ub1 = -3.191651871e-18 lub1 = 5.270333168e-25
+ uc1 = 3.615477057e-11 luc1 = -6.536546091e-18 puc1 = -7.346839693e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.87 nmos
* DC IV MOS Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.2025e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = 2.6e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 25000000.0
+ tnoib = 9900000.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {7.061484390e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -6.547863901e-08 wvth0 = -7.463212592e-09 pvth0 = 1.163888004e-15
+ k1 = 5.784727667e-01 lk1 = 1.758605004e-8
+ k2 = -6.613132729e-02 lk2 = -5.201017136e-09 wk2 = -2.444157735e-08 pk2 = 3.811663988e-15
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.851945716e+05 lvsat = -3.769572193e-03 wvsat = -1.512765376e-03 pvsat = 2.359157603e-10
+ ua = 3.111040417e-10 lua = -3.281278828e-16 wua = -5.426661083e-17 pua = 8.462877959e-24
+ ub = 2.545948883e-18 lub = 9.828143208e-27 wub = 1.331422922e-25 pub = -2.076354047e-32
+ uc = -3.661267122e-10 luc = 5.812183393e-17 wuc = 1.397863861e-16 puc = -2.179968692e-23
+ rdsw = 103.65
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = 6.517748496e-02 lu0 = -6.714810100e-09 wu0 = -2.708832491e-09 pu0 = 4.224424270e-16
+ a0 = 0.0
+ keta = -5.478114513e-01 lketa = 8.543119583e-08 wketa = 4.045286127e-07 pketa = -6.308623716e-14
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = 4.960995000e-01 lags = 9.408471298e-8
+ b0 = 0.0
+ b1 = 0.0
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.888714313e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 2.598017699e-08 wvoff = 4.817648731e-12 pvoff = -7.513123196e-19
+ nfactor = {-6.040426660e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 1.375221614e-06 wnfactor = 2.050968944e-06 pnfactor = -3.198486069e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = 2.553362249e-01 leta0 = -2.848513222e-8
+ etab = -1.545296712e-01 letab = 1.920177919e-8
+ dsub = 5.618342597e-01 ldsub = -3.801114066e-8
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 8.002976667e-02 lpclm = 3.604943839e-8
+ pdiblc1 = -3.995598333e+00 lpdiblc1 = 6.291956101e-07 wpdiblc1 = 4.235164736e-22 ppdiblc1 = -1.893266173e-29
+ pdiblc2 = 1.495856167e-02 lpdiblc2 = -4.078968419e-10
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 450000000.0
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.084666456e-03 lalpha0 = -5.583292809e-10 walpha0 = -7.342312099e-10 palpha0 = 1.145033572e-16
+ alpha1 = 0.0
+ beta0 = 1.566769616e+02 lbeta0 = -1.997416280e-05 wbeta0 = -4.364497377e-05 pbeta0 = 6.806433660e-12
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 1.4427e-15
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = -6.657438333e-02 lkt1 = -3.157763192e-8
+ kt2 = -7.388636000e-02 lkt2 = 6.851095592e-9
+ at = -1.179365980e+05 lat = 2.926660596e-02 wat = 6.171798645e-02 pat = -9.624919986e-9
+ ute = -1.816010500e+00 lute = 1.158872247e-8
+ ua1 = 2.281018004e-09 lua1 = -3.685532047e-16 wua1 = -6.456477888e-16 pua1 = 1.006887727e-22
+ ub1 = -4.854787000e-19 lub1 = 1.050056108e-25
+ uc1 = -1.097716290e-10 luc1 = 1.622067592e-17 wuc1 = -1.232595164e-32 puc1 = -7.346839693e-40
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 41000000.0
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.00275
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = 2.392894381e-10
+ cgso = 2.392894381e-10
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 2.310725e-11
+ cgdl = 2.310725e-11
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = 1.21071e-8
+ dwc = 2.6e-8
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0012094836
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = 3.230311424e-11
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = 1.795291232e-10
+ mjswgs = 0.8
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__nfet_01v8_lvt
