* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dlatn_1 D Q CLKN
X0 VDD a_n145_19 a_n78_109 VDD pmos_3p3 w=34 l=6
X1 a_n103_92 CLKN VDD VDD pmos_3p3 w=34 l=6
X2 Q a_n28_19 VDD VDD pmos_3p3 w=34 l=6
X3 VDD a_n135_14 a_n145_19 VDD pmos_3p3 w=34 l=6
X4 a_n112_109 D VDD VDD pmos_3p3 w=34 l=6
X5 a_n135_14 a_n103_92 a_n112_109 VDD pmos_3p3 w=34 l=6
X6 a_n78_19 a_n103_92 a_n135_14 GND nmos_3p3 w=17 l=6
X7 a_n103_92 CLKN GND GND nmos_3p3 w=17 l=6
X8 VDD a_n145_19 a_n28_19 VDD pmos_3p3 w=34 l=6
X9 a_n135_14 CLKN a_n109_19 GND nmos_3p3 w=17 l=6
X10 a_n109_19 D GND GND nmos_3p3 w=17 l=6
X11 GND a_n145_19 a_n78_19 GND nmos_3p3 w=17 l=6
X12 GND a_n135_14 a_n145_19 GND nmos_3p3 w=17 l=6
X13 a_n78_109 CLKN a_n135_14 VDD pmos_3p3 w=34 l=6
X14 GND a_n145_19 a_n28_19 GND nmos_3p3 w=17 l=6
X15 Q a_n28_19 GND GND nmos_3p3 w=17 l=6
.ends

