* NGSPICE file created from gf180mcu_osu_sc_9T_addf_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_9_70# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_110_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 S a_161_19# GND GND nmos_3p3 w=0.85u l=0.3u
X3 S a_161_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_195_19# B a_178_19# GND nmos_3p3 w=0.85u l=0.3u
X5 a_178_19# A a_161_19# GND nmos_3p3 w=0.85u l=0.3u
X6 a_195_70# B a_178_70# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_110_19# CI GND GND nmos_3p3 w=0.85u l=0.3u
X8 a_178_70# A a_161_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_59_19# CI a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X10 GND B a_110_19# GND nmos_3p3 w=0.85u l=0.3u
X11 a_110_70# CI VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 GND A a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X13 a_59_19# CI a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD B a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X15 CO a_59_19# GND GND nmos_3p3 w=0.85u l=0.3u
X16 VDD A a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X17 GND CI a_195_19# GND nmos_3p3 w=0.85u l=0.3u
X18 CO a_59_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 VDD CI a_195_70# VDD pmos_3p3 w=1.7u l=0.3u
X20 GND A a_76_19# GND nmos_3p3 w=0.85u l=0.3u
X21 a_161_19# a_59_19# a_110_19# GND nmos_3p3 w=0.85u l=0.3u
X22 a_76_19# B a_59_19# GND nmos_3p3 w=0.85u l=0.3u
X23 VDD A a_76_70# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_161_19# a_59_19# a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X25 a_9_19# B GND GND nmos_3p3 w=0.85u l=0.3u
X26 a_110_19# A GND GND nmos_3p3 w=0.85u l=0.3u
X27 a_76_70# B a_59_19# VDD pmos_3p3 w=1.7u l=0.3u
