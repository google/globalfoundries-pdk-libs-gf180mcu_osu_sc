# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__and2_1 0 0 ;
  SIZE 4.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.1 6.15 ;
        RECT 2.25 3.5 2.7 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.1 0.6 ;
        RECT 2.1 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.2 1.1 2.5 ;
        RECT 0.65 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.8 2.45 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 3.5 3.8 3.8 ;
        RECT 3.3 3.45 3.7 3.85 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 3.3 3.45 3.8 3.85 ;
      LAYER VIA12 ;
        RECT 3.42 3.52 3.68 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.45 1.65 5.2 ;
      RECT 2.75 2.1 3.05 2.6 ;
      RECT 1.4 2.2 3.05 2.5 ;
      RECT 0.7 1.45 1.65 1.7 ;
      RECT 0.7 0.95 0.95 1.7 ;
  END
END gf180mcu_osu_sc_gp9t3v3__and2_1
