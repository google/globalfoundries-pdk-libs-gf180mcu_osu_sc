* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_addf_1 A B CI S CO
X0 a_9_70 B VDD VDD pmos_3p3 w=34 l=6
X1 a_110_70 A VDD VDD pmos_3p3 w=34 l=6
X2 S a_161_19 GND GND nmos_3p3 w=17 l=6
X3 S a_161_19 VDD VDD pmos_3p3 w=34 l=6
X4 a_195_19 B a_178_19 GND nmos_3p3 w=17 l=6
X5 a_178_19 A a_161_19 GND nmos_3p3 w=17 l=6
X6 a_195_70 B a_178_70 VDD pmos_3p3 w=34 l=6
X7 a_110_19 CI GND GND nmos_3p3 w=17 l=6
X8 a_178_70 A a_161_19 VDD pmos_3p3 w=34 l=6
X9 a_59_19 CI a_9_19 GND nmos_3p3 w=17 l=6
X10 GND B a_110_19 GND nmos_3p3 w=17 l=6
X11 a_110_70 CI VDD VDD pmos_3p3 w=34 l=6
X12 GND A a_9_19 GND nmos_3p3 w=17 l=6
X13 a_59_19 CI a_9_70 VDD pmos_3p3 w=34 l=6
X14 VDD B a_110_70 VDD pmos_3p3 w=34 l=6
X15 CO a_59_19 GND GND nmos_3p3 w=17 l=6
X16 VDD A a_9_70 VDD pmos_3p3 w=34 l=6
X17 GND CI a_195_19 GND nmos_3p3 w=17 l=6
X18 CO a_59_19 VDD VDD pmos_3p3 w=34 l=6
X19 VDD CI a_195_70 VDD pmos_3p3 w=34 l=6
X20 GND A a_76_19 GND nmos_3p3 w=17 l=6
X21 a_161_19 a_59_19 a_110_19 GND nmos_3p3 w=17 l=6
X22 a_76_19 B a_59_19 GND nmos_3p3 w=17 l=6
X23 VDD A a_76_70 VDD pmos_3p3 w=34 l=6
X24 a_161_19 a_59_19 a_110_70 VDD pmos_3p3 w=34 l=6
X25 a_9_19 B GND GND nmos_3p3 w=17 l=6
X26 a_110_19 A GND GND nmos_3p3 w=17 l=6
X27 a_76_70 B a_59_19 VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
