magic
tech gf180mcuC
timestamp 1660079425
<< nwell >>
rect 0 97 32 159
<< metal1 >>
rect 0 147 32 159
rect 0 -3 32 9
<< labels >>
rlabel metal1 10 153 10 153 1 VDD
rlabel metal1 6 3 6 3 1 GND
<< end >>
