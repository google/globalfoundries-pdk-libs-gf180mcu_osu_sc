magic
tech gf180mcuC
timestamp 1659975287
<< nwell >>
rect 0 97 259 159
<< nmos >>
rect 19 16 25 33
rect 36 16 42 33
rect 52 16 58 33
rect 69 16 75 33
rect 80 16 86 33
rect 97 16 103 33
rect 108 16 114 33
rect 125 16 131 33
rect 136 16 142 33
rect 153 16 159 33
rect 185 16 191 33
rect 217 16 223 33
rect 234 16 240 33
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 52 106 58 140
rect 69 106 75 140
rect 80 106 86 140
rect 97 106 103 140
rect 108 106 114 140
rect 125 106 131 140
rect 136 106 142 140
rect 153 106 159 140
rect 185 106 191 140
rect 217 106 223 140
rect 234 106 240 140
<< ndiff >>
rect 9 31 19 33
rect 9 18 11 31
rect 16 18 19 31
rect 9 16 19 18
rect 25 31 36 33
rect 25 18 28 31
rect 33 18 36 31
rect 25 16 36 18
rect 42 16 52 33
rect 58 31 69 33
rect 58 18 61 31
rect 66 18 69 31
rect 58 16 69 18
rect 75 16 80 33
rect 86 23 97 33
rect 86 18 89 23
rect 94 18 97 23
rect 86 16 97 18
rect 103 16 108 33
rect 114 31 125 33
rect 114 18 117 31
rect 122 18 125 31
rect 114 16 125 18
rect 131 16 136 33
rect 142 31 153 33
rect 142 18 145 31
rect 150 18 153 31
rect 142 16 153 18
rect 159 31 169 33
rect 159 18 162 31
rect 167 18 169 31
rect 159 16 169 18
rect 175 24 185 33
rect 175 18 177 24
rect 182 18 185 24
rect 175 16 185 18
rect 191 31 201 33
rect 191 18 194 31
rect 199 18 201 31
rect 191 16 201 18
rect 207 31 217 33
rect 207 18 209 31
rect 214 18 217 31
rect 207 16 217 18
rect 223 31 234 33
rect 223 18 226 31
rect 231 18 234 31
rect 223 16 234 18
rect 240 31 250 33
rect 240 18 243 31
rect 248 18 250 31
rect 240 16 250 18
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 108 28 138
rect 33 108 36 138
rect 25 106 36 108
rect 42 106 52 140
rect 58 138 69 140
rect 58 108 61 138
rect 66 108 69 138
rect 58 106 69 108
rect 75 106 80 140
rect 86 138 97 140
rect 86 108 89 138
rect 94 108 97 138
rect 86 106 97 108
rect 103 106 108 140
rect 114 138 125 140
rect 114 123 117 138
rect 122 123 125 138
rect 114 106 125 123
rect 131 106 136 140
rect 142 138 153 140
rect 142 123 145 138
rect 150 123 153 138
rect 142 106 153 123
rect 159 138 169 140
rect 159 108 162 138
rect 167 108 169 138
rect 159 106 169 108
rect 175 138 185 140
rect 175 108 177 138
rect 182 108 185 138
rect 175 106 185 108
rect 191 138 201 140
rect 191 108 194 138
rect 199 108 201 138
rect 191 106 201 108
rect 207 138 217 140
rect 207 108 209 138
rect 214 108 217 138
rect 207 106 217 108
rect 223 138 234 140
rect 223 108 226 138
rect 231 108 234 138
rect 223 106 234 108
rect 240 138 250 140
rect 240 108 243 138
rect 248 108 250 138
rect 240 106 250 108
<< ndiffc >>
rect 11 18 16 31
rect 28 18 33 31
rect 61 18 66 31
rect 89 18 94 23
rect 117 18 122 31
rect 145 18 150 31
rect 162 18 167 31
rect 177 18 182 24
rect 194 18 199 31
rect 209 18 214 31
rect 226 18 231 31
rect 243 18 248 31
<< pdiffc >>
rect 11 108 16 138
rect 28 108 33 138
rect 61 108 66 138
rect 89 108 94 138
rect 117 123 122 138
rect 145 123 150 138
rect 162 108 167 138
rect 177 108 182 138
rect 194 108 199 138
rect 209 108 214 138
rect 226 108 231 138
rect 243 108 248 138
<< psubdiff >>
rect 9 7 18 9
rect 9 2 11 7
rect 16 2 18 7
rect 9 0 18 2
rect 33 7 42 9
rect 33 2 35 7
rect 40 2 42 7
rect 33 0 42 2
rect 57 7 66 9
rect 57 2 59 7
rect 64 2 66 7
rect 57 0 66 2
rect 81 7 90 9
rect 81 2 83 7
rect 88 2 90 7
rect 81 0 90 2
rect 105 7 114 9
rect 105 2 107 7
rect 112 2 114 7
rect 105 0 114 2
rect 129 7 138 9
rect 129 2 131 7
rect 136 2 138 7
rect 129 0 138 2
rect 153 7 162 9
rect 153 2 155 7
rect 160 2 162 7
rect 153 0 162 2
rect 177 7 186 9
rect 177 2 179 7
rect 184 2 186 7
rect 177 0 186 2
rect 201 7 210 9
rect 201 2 203 7
rect 208 2 210 7
rect 201 0 210 2
rect 225 7 234 9
rect 225 2 227 7
rect 232 2 234 7
rect 225 0 234 2
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
rect 81 154 90 156
rect 81 149 83 154
rect 88 149 90 154
rect 81 147 90 149
rect 105 154 114 156
rect 105 149 107 154
rect 112 149 114 154
rect 105 147 114 149
rect 129 154 138 156
rect 129 149 131 154
rect 136 149 138 154
rect 129 147 138 149
rect 153 154 162 156
rect 153 149 155 154
rect 160 149 162 154
rect 153 147 162 149
rect 177 154 186 156
rect 177 149 179 154
rect 184 149 186 154
rect 177 147 186 149
rect 201 154 210 156
rect 201 149 203 154
rect 208 149 210 154
rect 201 147 210 149
rect 225 154 234 156
rect 225 149 227 154
rect 232 149 234 154
rect 225 147 234 149
<< psubdiffcont >>
rect 11 2 16 7
rect 35 2 40 7
rect 59 2 64 7
rect 83 2 88 7
rect 107 2 112 7
rect 131 2 136 7
rect 155 2 160 7
rect 179 2 184 7
rect 203 2 208 7
rect 227 2 232 7
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
rect 83 149 88 154
rect 107 149 112 154
rect 131 149 136 154
rect 155 149 160 154
rect 179 149 184 154
rect 203 149 208 154
rect 227 149 232 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 52 140 58 145
rect 69 140 75 145
rect 80 140 86 145
rect 97 140 103 145
rect 108 140 114 145
rect 125 140 131 145
rect 136 140 142 145
rect 153 140 159 145
rect 185 140 191 145
rect 217 140 223 145
rect 234 140 240 145
rect 19 88 25 106
rect 19 86 31 88
rect 19 80 23 86
rect 29 80 31 86
rect 19 78 31 80
rect 19 33 25 78
rect 36 75 42 106
rect 52 88 58 106
rect 52 86 62 88
rect 52 80 54 86
rect 60 80 62 86
rect 52 78 62 80
rect 36 73 48 75
rect 36 67 40 73
rect 46 67 48 73
rect 36 65 48 67
rect 36 33 42 65
rect 69 61 75 106
rect 80 101 86 106
rect 97 101 103 106
rect 80 99 103 101
rect 80 94 83 99
rect 81 93 83 94
rect 89 94 103 99
rect 89 93 91 94
rect 81 89 91 93
rect 108 61 114 106
rect 125 88 131 106
rect 121 86 131 88
rect 121 80 123 86
rect 129 80 131 86
rect 121 78 131 80
rect 136 75 142 106
rect 153 88 159 106
rect 153 86 163 88
rect 153 80 155 86
rect 161 80 163 86
rect 153 78 163 80
rect 135 73 145 75
rect 135 67 137 73
rect 143 67 145 73
rect 135 65 145 67
rect 121 61 131 62
rect 52 60 131 61
rect 52 55 123 60
rect 52 33 58 55
rect 121 54 123 55
rect 129 54 131 60
rect 121 52 131 54
rect 65 47 75 49
rect 81 47 91 49
rect 65 41 67 47
rect 73 41 75 47
rect 65 39 75 41
rect 69 33 75 39
rect 80 41 83 47
rect 89 41 103 47
rect 80 39 103 41
rect 80 33 86 39
rect 97 33 103 39
rect 108 46 118 48
rect 108 40 110 46
rect 116 40 118 46
rect 108 38 118 40
rect 108 33 114 38
rect 125 33 131 52
rect 136 33 142 65
rect 153 33 159 78
rect 185 62 191 106
rect 217 62 223 106
rect 234 88 240 106
rect 228 86 240 88
rect 228 80 230 86
rect 236 80 240 86
rect 228 78 240 80
rect 179 60 191 62
rect 179 54 181 60
rect 187 54 191 60
rect 179 52 191 54
rect 211 60 223 62
rect 211 54 215 60
rect 221 54 223 60
rect 211 52 223 54
rect 185 33 191 52
rect 217 33 223 52
rect 234 33 240 78
rect 19 11 25 16
rect 36 11 42 16
rect 52 11 58 16
rect 69 11 75 16
rect 80 11 86 16
rect 97 11 103 16
rect 108 11 114 16
rect 125 11 131 16
rect 136 11 142 16
rect 153 11 159 16
rect 185 11 191 16
rect 217 11 223 16
rect 234 11 240 16
<< polycontact >>
rect 23 80 29 86
rect 54 80 60 86
rect 40 67 46 73
rect 83 93 89 99
rect 123 80 129 86
rect 155 80 161 86
rect 137 67 143 73
rect 123 54 129 60
rect 67 41 73 47
rect 83 41 89 47
rect 110 40 116 46
rect 230 80 236 86
rect 181 54 187 60
rect 215 54 221 60
<< metal1 >>
rect 0 154 259 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 83 154
rect 89 148 107 154
rect 113 148 131 154
rect 137 148 155 154
rect 161 148 179 154
rect 185 148 203 154
rect 209 148 227 154
rect 233 148 259 154
rect 0 147 259 148
rect 11 138 16 140
rect 11 49 16 108
rect 28 138 33 147
rect 28 106 33 108
rect 61 138 66 140
rect 61 101 66 108
rect 89 138 94 147
rect 117 138 122 140
rect 117 121 122 123
rect 145 138 150 147
rect 145 121 150 123
rect 162 138 167 140
rect 89 106 94 108
rect 99 116 122 121
rect 28 96 66 101
rect 28 86 33 96
rect 81 93 83 99
rect 89 93 91 99
rect 21 80 23 86
rect 29 80 33 86
rect 52 80 54 86
rect 60 80 67 86
rect 73 80 75 86
rect 10 47 16 49
rect 28 47 33 80
rect 38 67 40 73
rect 46 67 48 73
rect 67 47 73 80
rect 83 47 89 93
rect 99 71 104 116
rect 134 93 136 99
rect 142 93 144 99
rect 162 97 167 108
rect 177 138 182 147
rect 177 106 182 108
rect 194 138 199 140
rect 98 66 104 71
rect 110 80 123 86
rect 129 80 131 86
rect 28 42 48 47
rect 10 39 16 41
rect 11 31 16 39
rect 40 33 48 42
rect 65 41 67 47
rect 73 41 75 47
rect 81 41 83 47
rect 89 41 91 47
rect 98 34 103 66
rect 110 46 116 80
rect 136 73 142 93
rect 162 92 178 97
rect 153 80 155 86
rect 161 80 163 86
rect 172 73 178 92
rect 135 67 137 73
rect 143 67 145 73
rect 162 68 178 73
rect 162 60 168 68
rect 181 60 187 62
rect 194 60 199 108
rect 209 138 214 140
rect 209 86 214 108
rect 226 138 231 147
rect 226 106 231 108
rect 243 138 248 140
rect 243 100 248 108
rect 243 99 253 100
rect 243 93 245 99
rect 251 93 253 99
rect 243 92 252 93
rect 209 80 230 86
rect 236 80 238 86
rect 121 54 123 60
rect 129 54 131 60
rect 179 54 181 60
rect 187 54 189 60
rect 194 54 215 60
rect 221 54 223 60
rect 162 52 168 54
rect 108 40 110 46
rect 116 40 118 46
rect 11 16 16 18
rect 28 31 33 33
rect 40 31 66 33
rect 40 28 61 31
rect 28 9 33 18
rect 98 29 117 34
rect 123 28 125 34
rect 145 31 150 33
rect 61 16 66 18
rect 89 23 94 25
rect 89 9 94 18
rect 117 16 122 18
rect 145 9 150 18
rect 162 31 167 52
rect 181 37 187 54
rect 179 31 181 37
rect 187 31 189 37
rect 194 31 199 54
rect 231 43 236 80
rect 162 16 167 18
rect 177 24 182 26
rect 177 9 182 18
rect 194 16 199 18
rect 209 38 236 43
rect 209 31 214 38
rect 209 16 214 18
rect 226 31 231 33
rect 226 9 231 18
rect 243 31 248 92
rect 243 16 248 18
rect 0 8 259 9
rect 0 2 11 8
rect 17 2 35 8
rect 41 2 59 8
rect 65 2 83 8
rect 89 2 107 8
rect 113 2 131 8
rect 137 2 155 8
rect 161 2 179 8
rect 185 2 203 8
rect 209 2 227 8
rect 233 2 259 8
rect 0 -3 259 2
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 83 149 88 154
rect 88 149 89 154
rect 83 148 89 149
rect 107 149 112 154
rect 112 149 113 154
rect 107 148 113 149
rect 131 149 136 154
rect 136 149 137 154
rect 131 148 137 149
rect 155 149 160 154
rect 160 149 161 154
rect 155 148 161 149
rect 179 149 184 154
rect 184 149 185 154
rect 179 148 185 149
rect 203 149 208 154
rect 208 149 209 154
rect 203 148 209 149
rect 227 149 232 154
rect 232 149 233 154
rect 227 148 233 149
rect 67 80 73 86
rect 10 41 16 47
rect 40 67 46 73
rect 136 93 142 99
rect 123 80 129 86
rect 83 41 89 47
rect 155 80 161 86
rect 137 67 143 73
rect 245 93 251 99
rect 230 80 236 86
rect 123 54 129 60
rect 162 54 168 60
rect 215 54 221 60
rect 117 31 123 34
rect 117 28 122 31
rect 122 28 123 31
rect 181 31 187 37
rect 11 7 17 8
rect 11 2 16 7
rect 16 2 17 7
rect 35 7 41 8
rect 35 2 40 7
rect 40 2 41 7
rect 59 7 65 8
rect 59 2 64 7
rect 64 2 65 7
rect 83 7 89 8
rect 83 2 88 7
rect 88 2 89 7
rect 107 7 113 8
rect 107 2 112 7
rect 112 2 113 7
rect 131 7 137 8
rect 131 2 136 7
rect 136 2 137 7
rect 155 7 161 8
rect 155 2 160 7
rect 160 2 161 7
rect 179 7 185 8
rect 179 2 184 7
rect 184 2 185 7
rect 203 7 209 8
rect 203 2 208 7
rect 208 2 209 7
rect 227 7 233 8
rect 227 2 232 7
rect 232 2 233 7
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 130 154 138 155
rect 154 154 162 155
rect 178 154 186 155
rect 202 154 210 155
rect 226 154 234 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 81 148 83 154
rect 89 148 91 154
rect 105 148 107 154
rect 113 148 115 154
rect 129 148 131 154
rect 137 148 139 154
rect 153 148 155 154
rect 161 148 163 154
rect 177 148 179 154
rect 185 148 187 154
rect 201 148 203 154
rect 209 148 211 154
rect 225 148 227 154
rect 233 148 235 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 130 147 138 148
rect 154 147 162 148
rect 178 147 186 148
rect 202 147 210 148
rect 226 147 234 148
rect 135 99 143 100
rect 244 99 252 100
rect 134 93 136 99
rect 142 93 198 99
rect 243 93 245 99
rect 251 93 253 99
rect 135 92 143 93
rect 65 86 74 87
rect 121 86 131 87
rect 154 86 162 87
rect 65 80 67 86
rect 73 80 123 86
rect 129 80 155 86
rect 161 80 163 86
rect 65 79 74 80
rect 121 79 131 80
rect 154 79 162 80
rect 38 73 48 74
rect 136 73 144 74
rect 35 67 40 73
rect 46 67 51 73
rect 135 67 137 73
rect 143 67 145 73
rect 38 66 48 67
rect 136 66 144 67
rect 122 60 130 61
rect 161 60 169 61
rect 192 60 198 93
rect 244 92 252 93
rect 229 86 237 87
rect 228 80 230 86
rect 236 80 238 86
rect 229 79 237 80
rect 214 60 222 61
rect 121 54 123 60
rect 129 54 162 60
rect 168 54 171 60
rect 192 54 215 60
rect 221 54 223 60
rect 122 53 130 54
rect 161 53 169 54
rect 214 53 222 54
rect 9 47 17 48
rect 82 47 90 48
rect 8 41 10 47
rect 16 41 83 47
rect 89 41 91 47
rect 9 40 17 41
rect 82 40 90 41
rect 180 37 188 38
rect 116 34 124 35
rect 170 34 181 37
rect 115 28 117 34
rect 123 31 181 34
rect 187 31 189 37
rect 123 30 188 31
rect 123 28 176 30
rect 116 27 124 28
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 82 8 90 9
rect 106 8 114 9
rect 130 8 138 9
rect 154 8 162 9
rect 178 8 186 9
rect 202 8 210 9
rect 226 8 234 9
rect 9 2 11 8
rect 17 2 19 8
rect 33 2 35 8
rect 41 2 43 8
rect 57 2 59 8
rect 65 2 67 8
rect 81 2 83 8
rect 89 2 91 8
rect 105 2 107 8
rect 113 2 115 8
rect 129 2 131 8
rect 137 2 139 8
rect 153 2 155 8
rect 161 2 163 8
rect 177 2 179 8
rect 185 2 187 8
rect 201 2 203 8
rect 209 2 211 8
rect 225 2 227 8
rect 233 2 235 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
rect 82 1 90 2
rect 106 1 114 2
rect 130 1 138 2
rect 154 1 162 2
rect 178 1 186 2
rect 202 1 210 2
rect 226 1 234 2
<< labels >>
rlabel metal2 248 96 248 96 1 Q
port 4 n
rlabel metal2 43 70 43 70 1 D
port 1 n
rlabel metal2 13 5 13 5 1 GND
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 233 83 233 83 1 QN
port 6 n
rlabel metal2 158 83 158 83 1 CLKN
port 7 n
<< end >>
