* NGSPICE file created from gf180mcu_osu_sc_9T_dffn_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_42_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_125_19# a_53_38# a_114_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_86_70# a_53_38# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD a_161_42# a_148_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 GND a_9_19# a_86_19# GND nmos_3p3 w=0.85u l=0.3u
X5 a_19_14# a_53_38# a_42_19# GND nmos_3p3 w=0.85u l=0.3u
X6 GND a_161_42# QN GND nmos_3p3 w=0.85u l=0.3u
X7 VDD a_9_19# a_86_70# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_19_14# CLKN a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X9 VDD a_161_42# QN VDD pmos_3p3 w=1.7u l=0.3u
X10 GND a_19_14# a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X11 a_53_38# CLKN GND GND nmos_3p3 w=0.85u l=0.3u
X12 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X13 a_53_38# CLKN VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 a_148_19# a_53_38# a_125_19# GND nmos_3p3 w=0.85u l=0.3u
X15 Q QN GND GND nmos_3p3 w=0.85u l=0.3u
X16 a_114_19# a_9_19# GND GND nmos_3p3 w=0.85u l=0.3u
X17 a_161_42# a_125_19# GND GND nmos_3p3 w=0.85u l=0.3u
X18 a_148_70# CLKN a_125_19# VDD pmos_3p3 w=1.7u l=0.3u
X19 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X20 a_114_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X21 a_161_42# a_125_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 a_42_19# D GND GND nmos_3p3 w=0.85u l=0.3u
X23 a_125_19# CLKN a_114_19# GND nmos_3p3 w=0.85u l=0.3u
X24 a_86_19# CLKN a_19_14# GND nmos_3p3 w=0.85u l=0.3u
X25 GND a_161_42# a_148_19# GND nmos_3p3 w=0.85u l=0.3u
