* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsn_1 D Q QN CLK SN VDD VSS
X0 a_75_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_147_21# a_242_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_242_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VSS SN a_108_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS CLK a_85_83# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_85_16# a_85_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_85_16# a_85_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_75_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X8 VDD a_168_70# a_164_111# VDD pfet_03p3 w=1.7u l=0.3u
X9 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VDD SN SN VDD pfet_03p3 w=1.7u l=0.3u
X11 SN a_34_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X12 a_147_21# a_85_16# a_136_111# VDD pfet_03p3 w=1.7u l=0.3u
X13 a_164_111# a_85_83# a_147_21# VDD pfet_03p3 w=1.7u l=0.3u
X14 VDD CLK a_85_83# VDD pfet_03p3 w=1.7u l=0.3u
X15 a_261_21# a_147_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 VSS a_168_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X17 a_136_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X18 VDD SN a_108_111# VDD pfet_03p3 w=1.7u l=0.3u
X19 a_136_21# SN VSS VSS nfet_03p3 w=0.85u l=0.3u
X20 a_164_21# a_85_16# a_147_21# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_168_70# SN a_261_21# VSS nfet_03p3 w=0.85u l=0.3u
X22 a_108_111# a_85_16# a_34_16# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_147_21# a_85_83# a_136_21# VSS nfet_03p3 w=0.85u l=0.3u
X24 VSS a_168_70# a_164_21# VSS nfet_03p3 w=0.85u l=0.3u
X25 a_34_16# a_85_83# a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_29_21# SN SN VSS nfet_03p3 w=0.85u l=0.3u
X27 a_34_16# a_85_16# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X28 VDD a_168_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X29 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 VSS a_34_16# a_29_21# VSS nfet_03p3 w=0.85u l=0.3u
X31 a_108_21# a_85_83# a_34_16# VSS nfet_03p3 w=0.85u l=0.3u
.ends
