* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.subckt  sky130_fd_pr__esd_nfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__esd_nfet_g5v0d10v5.0 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.7495e-05 wmax = 1.7505e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_0}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_0}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109000+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_0}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_0}
+ ub = {1.4129e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_0}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_0}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_0}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_0}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_0}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_0}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_0}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_0}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_0}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_0}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_0}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_0}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_0}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_0}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_0}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.1 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 1.9495e-05 wmax = 1.9505e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_1}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_1}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109850+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_1}
+ ua = {1.6364e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_1}
+ ub = {1.0455e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_1}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_1}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_1}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_1}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_1}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_1}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_1}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_1}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_1}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_1}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_1}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_1}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_1}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_1}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_1}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.2 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.1495e-05 wmax = 2.1505e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_2}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_2}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {107440+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_2}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_2}
+ ub = {1.4129e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_2}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_2}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_2}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_2}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_2}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_2}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_2}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_2}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_2}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_2}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_2}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_2}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_2}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_2}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_2}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.3 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.3495e-05 wmax = 2.3505e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_3}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_3}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108170+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_3}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_3}
+ ub = {1.4129e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_3}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_3}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_3}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_3}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_3}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_3}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_3}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_3}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_3}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_3}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_3}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_3}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_3}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_3}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_3}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.4 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 2.6495e-05 wmax = 2.6505e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_4}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_4}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108170+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_4}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_4}
+ ub = {1.5358e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_4}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_4}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_4}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_4}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_4}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_4}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_4}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_4}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_4}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_4}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_4}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_4}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_4}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_4}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_4}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.5 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 3.0245e-05 wmax = 3.0255e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.798+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_5}
+ k1 = 0.76281
+ k2 = {-0.071923+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_5}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {89500+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_5}
+ ua = {1.0364e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_5}
+ ub = {1.5358e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_5}
+ uc = 5.215e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_5}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.060184+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_5}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_5}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_5}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_5}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_5}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_5}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_5}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_5}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_5}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_5}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_5}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_5}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_5}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.6 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 3.0245e-05 wmax = 3.0255e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.814+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_6}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_6}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108170+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_6}
+ ua = {1.3637e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_6}
+ ub = {1.5358e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_6}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_6}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_6}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_6}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_6}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_6}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_6}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_6}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_6}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_6}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_6}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_6}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_6}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_6}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_6}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.7 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 4.0305e-05 wmax = 4.0315e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.805+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_7}
+ k1 = 0.76281
+ k2 = {-0.081731+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_7}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108170+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_7}
+ ua = {1.1962e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_7}
+ ub = {1.8283e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_7}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_7}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.066871+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_7}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_7}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_7}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_7}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_7}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_7}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_7}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_7}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_7}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 5.088e+8
+ pscbe2 = 2.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.6845e-5
+ alpha1 = 0.37039
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_7}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_7}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_7}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_7}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.8 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 5.0985e-05 wmax = 5.0995e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.807+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_8}
+ k1 = 0.75481
+ k2 = {-0.033568+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_8}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {91046+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_8}
+ ua = {1.1962e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_8}
+ ub = {1.7552e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_8}
+ uc = 8.4519e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_8}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.064299+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_8}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_8}
+ keta = {-0.041308+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_8}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_8}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_8}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_8}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_8}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_8}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_8}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0018
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 4.2400001e+9
+ pscbe2 = 1.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 4.9691e-5
+ alpha1 = 0.8052
+ beta0 = 38.234
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_8}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_8}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_8}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_8}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.9 nmos
* DC IV MOS Parameters
+ lmin = 5.45e-07 lmax = 5.55e-07 wmin = 5.0985e-05 wmax = 5.0995e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.815+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_9}
+ k1 = 0.76281
+ k2 = {-0.072974+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_9}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109170+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_9}
+ ua = {1.1962e-009+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_9}
+ ub = {1.8283e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_9}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_9}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.064299+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_9}
+ a0 = {0.1054+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_9}
+ keta = {-0.057372+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.48+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_9}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_9}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_9}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_9}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_9}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.21835+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_9}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_9}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 4.2400001e+9
+ pscbe2 = 1.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 2.8558e-5
+ alpha1 = 0.8052
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_9}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_9}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_9}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_9}
+ kt2 = -0.015814
+ at = 38574.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 4.7889e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.model sky130_fd_pr__esd_nfet_g5v0d10v5.10 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 5.395e-06 wmax = 5.405e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {3.6e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {-5.8413e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = 0.0
+ dwb = 3.3727471e-12
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.577
+ rnoib = 0.5164
+ tnoia = 1.5
+ tnoib = 3.5
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__esd_nfet_g5v0d10v5__toxe_mult}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__esd_nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82+sky130_fd_pr__esd_nfet_g5v0d10v5__vth0_diff_10}
+ k1 = 0.76281
+ k2 = {-0.061842+sky130_fd_pr__esd_nfet_g5v0d10v5__k2_diff_10}
+ k3 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.5
+ dvt2 = -0.001152
+ dvt0w = 0.0
+ dvt1w = 5215200.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108590+sky130_fd_pr__esd_nfet_g5v0d10v5__vsat_diff_10}
+ ua = {6e-010+sky130_fd_pr__esd_nfet_g5v0d10v5__ua_diff_10}
+ ub = {1.6038e-018+sky130_fd_pr__esd_nfet_g5v0d10v5__ub_diff_10}
+ uc = 4.4957e-11
+ rdsw = {566.95+sky130_fd_pr__esd_nfet_g5v0d10v5__rdsw_diff_10}
+ prwb = 0.015804
+ prwg = 5.4e-13
+ wr = 1.0
+ u0 = {0.057246+sky130_fd_pr__esd_nfet_g5v0d10v5__u0_diff_10}
+ a0 = {0.00+sky130_fd_pr__esd_nfet_g5v0d10v5__a0_diff_10}
+ keta = {-0.045533+sky130_fd_pr__esd_nfet_g5v0d10v5__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {1+sky130_fd_pr__esd_nfet_g5v0d10v5__ags_diff_10}
+ b0 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b0_diff_10}
+ b1 = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__voff_diff_10}
+ nfactor = {0.114+sky130_fd_pr__esd_nfet_g5v0d10v5__nfactor_diff_10}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__tvoff_diff_10}
+ cit = -0.0007128
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.0e-12
+ eta0 = {0.059173+sky130_fd_pr__esd_nfet_g5v0d10v5__eta0_diff_10}
+ etab = -0.0031079
+ dsub = 0.5
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23915+sky130_fd_pr__esd_nfet_g5v0d10v5__pclm_diff_10}
+ pdiblc1 = 0.09332
+ pdiblc2 = 0.0
+ pdiblcb = -0.26831
+ drout = 0.2822
+ pscbe1 = 4.2400001e+9
+ pscbe2 = 1.0e-8
+ pvag = 1.9901676
+ delta = 0.0445
+ alpha0 = 4.6061e-5
+ alpha1 = 0.8052
+ beta0 = 39.827
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.4829e-007+sky130_fd_pr__esd_nfet_g5v0d10v5__agidl_diff_10}
+ bgidl = {2.4214e+009+sky130_fd_pr__esd_nfet_g5v0d10v5__bgidl_diff_10}
+ cgidl = {10120+sky130_fd_pr__esd_nfet_g5v0d10v5__cgidl_diff_10}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.34313+sky130_fd_pr__esd_nfet_g5v0d10v5__kt1_diff_10}
+ kt2 = -0.015814289
+ at = 30614.0
+ ute = -1.4571
+ ua1 = 3.4582e-9
+ ub1 = -3.4538e-18
+ uc1 = 1.6097e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 2.0
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__esd_nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__esd_nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__esd_nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__esd_nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
.ends sky130_fd_pr__esd_nfet_g5v0d10v5
