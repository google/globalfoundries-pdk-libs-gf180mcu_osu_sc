# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi21_1 0 0 ;
  SIZE 3.9 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 3.9 6.35 ;
        RECT 1.4 4.35 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 2.95 0 3.2 1.5 ;
        RECT 0.7 0 0.95 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 2.95 2.1 3.25 ;
      LAYER Metal2 ;
        RECT 1.6 2.9 2.1 3.3 ;
      LAYER Via1 ;
        RECT 1.72 2.97 1.98 3.23 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.35 2.3 2.85 2.6 ;
      LAYER Metal2 ;
        RECT 2.35 2.25 2.85 2.65 ;
      LAYER Via1 ;
        RECT 2.47 2.32 2.73 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 3.6 3.5 3.9 ;
        RECT 3.1 1.75 3.35 5.3 ;
        RECT 2.1 1.75 3.35 2 ;
        RECT 2.1 1.05 2.35 2 ;
      LAYER Metal2 ;
        RECT 3 3.55 3.5 3.95 ;
      LAYER Via1 ;
        RECT 3.12 3.62 3.38 3.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 2.25 3.85 2.5 5.3 ;
      RECT 0.55 3.85 0.8 5.3 ;
      RECT 0.55 3.85 2.5 4.1 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi21_1
