# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__mux2_1 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 3.45 2.85 3.85 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.75 4.1 4.25 4.5 ;
        RECT 3.95 0.95 4.2 7.15 ;
      LAYER MET2 ;
        RECT 3.75 4.1 4.25 4.5 ;
      LAYER VIA12 ;
        RECT 3.87 4.17 4.13 4.43 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.85 1.05 3.15 ;
      LAYER MET2 ;
        RECT 0.55 2.8 1.05 3.2 ;
      LAYER VIA12 ;
        RECT 0.67 2.87 0.93 3.13 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.75 3.5 5.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
      LAYER MET2 ;
        RECT 3 4.75 3.5 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 4.82 3.38 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.4 4.15 2 4.45 ;
      RECT 1.4 2.2 2 2.5 ;
  END
END gf180mcu_osu_sc_gp12t3v3__mux2_1
