# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_8 0 0 ;
  SIZE 9.05 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 9.05 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.05 0.6 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 3.5 7.75 3.8 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 2.25 2.95 7.6 3.25 ;
        RECT 2.25 2.05 7.6 2.35 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 7.25 3.45 7.75 3.85 ;
      LAYER VIA12 ;
        RECT 7.37 3.52 7.63 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_8
