# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_oai21_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_oai21_1 0 -0.15 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.35 0.95 3.65 ;
      LAYER MET2 ;
        RECT 0.45 3.3 0.95 3.7 ;
      LAYER VIA12 ;
        RECT 0.57 3.37 0.83 3.63 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4 1.95 4.3 ;
      LAYER MET2 ;
        RECT 1.45 3.95 1.95 4.35 ;
      LAYER VIA12 ;
        RECT 1.57 4.02 1.83 4.28 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 3.35 2.7 3.65 ;
      LAYER MET2 ;
        RECT 2.2 3.3 2.7 3.7 ;
      LAYER VIA12 ;
        RECT 2.32 3.37 2.58 3.63 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 3.9 7.95 ;
        RECT 2.95 5.3 3.2 7.95 ;
        RECT 0.65 5.3 0.9 7.95 ;
      LAYER MET2 ;
        RECT 2.85 7.4 3.35 7.7 ;
        RECT 2.9 7.35 3.3 7.75 ;
        RECT 1.65 7.4 2.15 7.7 ;
        RECT 1.7 7.35 2.1 7.75 ;
        RECT 0.45 7.4 0.95 7.7 ;
        RECT 0.5 7.35 0.9 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
        RECT 1.77 7.42 2.03 7.68 ;
        RECT 2.97 7.42 3.23 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 3.9 0.45 ;
        RECT 1.35 -0.15 1.6 1.35 ;
      LAYER MET2 ;
        RECT 2.85 0.1 3.35 0.4 ;
        RECT 2.9 0.05 3.3 0.45 ;
        RECT 1.65 0.1 2.15 0.4 ;
        RECT 1.7 0.05 2.1 0.45 ;
        RECT 0.45 0.1 0.95 0.4 ;
        RECT 0.5 0.05 0.9 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
        RECT 1.77 0.12 2.03 0.38 ;
        RECT 2.97 0.12 3.23 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 4.65 3.35 4.95 ;
        RECT 3.05 0.8 3.3 2.35 ;
        RECT 2.95 2.1 3.2 4.95 ;
        RECT 2.1 4.65 2.35 7 ;
      LAYER MET2 ;
        RECT 2.85 4.6 3.35 5 ;
      LAYER VIA12 ;
        RECT 2.97 4.67 3.23 4.93 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.6 2.45 1.85 ;
      RECT 2.2 0.8 2.45 1.85 ;
      RECT 0.5 0.8 0.75 1.85 ;
  END
END gf180mcu_osu_sc_12T_oai21_1
