* NGSPICE file created from gf180mcu_osu_sc_9T_buf_2.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 GND a_9_19# Y GND nmos_3p3 w=0.85u l=0.3u
X2 GND A a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X3 VDD a_9_19# Y VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 Y a_9_19# GND GND nmos_3p3 w=0.85u l=0.3u
