VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addf_1 0 0 ;
  SIZE 14 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 14 8.1 ;
        RECT 12.35 5.45 12.6 8.1 ;
        RECT 10.75 5.45 11 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14 0.6 ;
        RECT 12.35 0 12.6 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 6.5 0 6.75 1.45 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.7 3.5 9.2 3.8 ;
        RECT 4.6 3.5 5.1 3.8 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.5 9.2 3.8 ;
        RECT 8.75 3.45 9.15 3.85 ;
        RECT 4.65 3.45 5.05 3.85 ;
        RECT 0.65 3.45 1.05 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
        RECT 4.72 3.52 4.98 3.78 ;
        RECT 8.82 3.52 9.08 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.55 4.15 10.05 4.45 ;
        RECT 3.6 4.15 6.25 4.45 ;
        RECT 1.5 4.15 2 4.45 ;
      LAYER MET2 ;
        RECT 5.75 4.15 10.05 4.45 ;
        RECT 9.6 4.1 10 4.5 ;
        RECT 5.8 4.1 6.2 4.5 ;
        RECT 1.5 4.15 4.1 4.45 ;
        RECT 3.65 4.1 4.05 4.5 ;
        RECT 1.55 4.1 1.95 4.5 ;
      LAYER VIA12 ;
        RECT 1.62 4.17 1.88 4.43 ;
        RECT 3.72 4.17 3.98 4.43 ;
        RECT 5.87 4.17 6.13 4.43 ;
        RECT 9.67 4.17 9.93 4.43 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.05 2.2 10.55 2.5 ;
        RECT 6.65 2.2 7.15 2.5 ;
        RECT 2.35 2.85 2.85 3.15 ;
      LAYER MET2 ;
        RECT 2.45 2.2 10.55 2.5 ;
        RECT 10.1 2.15 10.5 2.55 ;
        RECT 10.15 2.1 10.45 2.55 ;
        RECT 6.7 2.15 7.1 2.55 ;
        RECT 6.75 2.1 7.05 2.55 ;
        RECT 2.35 2.85 2.85 3.15 ;
        RECT 2.4 2.8 2.8 3.2 ;
        RECT 2.45 2.2 2.75 3.2 ;
      LAYER VIA12 ;
        RECT 2.47 2.87 2.73 3.13 ;
        RECT 6.77 2.22 7.03 2.48 ;
        RECT 10.17 2.22 10.43 2.48 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.2 2.85 13.75 3.15 ;
        RECT 13.2 2.8 13.6 3.2 ;
        RECT 13.2 0.95 13.45 7.15 ;
      LAYER MET2 ;
        RECT 13.25 2.85 13.75 3.15 ;
        RECT 13.3 2.8 13.7 3.2 ;
      LAYER VIA12 ;
        RECT 13.37 2.87 13.63 3.13 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.6 4.15 12 4.45 ;
        RECT 11.6 0.95 11.85 7.15 ;
      LAYER MET2 ;
        RECT 11.5 4.15 12 4.45 ;
        RECT 11.55 4.1 11.95 4.5 ;
      LAYER VIA12 ;
        RECT 11.62 4.17 11.88 4.43 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 12.5 2.8 12.9 3.2 ;
      RECT 7.5 2.8 7.9 3.2 ;
      RECT 7.45 2.85 12.95 3.15 ;
      RECT 12.55 2.75 12.85 3.2 ;
    LAYER VIA12 ;
      RECT 12.57 2.87 12.83 3.13 ;
      RECT 7.57 2.87 7.83 3.13 ;
    LAYER MET1 ;
      RECT 8.2 0.95 8.45 7.15 ;
      RECT 8.2 2.85 11.35 3.15 ;
      RECT 3.1 0.95 3.35 7.15 ;
      RECT 3.1 2.85 7.95 3.15 ;
      RECT 5.65 1.7 7.6 1.95 ;
      RECT 7.35 0.95 7.6 1.95 ;
      RECT 5.65 0.95 5.9 1.95 ;
      RECT 7.35 4.95 7.6 7.15 ;
      RECT 5.65 4.95 5.9 7.15 ;
      RECT 5.65 4.95 7.6 5.2 ;
      RECT 0.55 2.05 2.5 2.3 ;
      RECT 2.25 0.95 2.5 2.3 ;
      RECT 0.55 0.95 0.8 2.3 ;
      RECT 2.25 4.95 2.5 7.15 ;
      RECT 0.55 4.95 0.8 7.15 ;
      RECT 0.55 4.95 2.5 5.2 ;
      RECT 12.45 2.85 12.95 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addf_1

MACRO gf180mcu_osu_sc_gp12t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addh_1 0 0 ;
  SIZE 8.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 8.1 8.1 ;
        RECT 6.4 5.45 6.65 8.1 ;
        RECT 3.85 5.45 4.1 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.1 0.6 ;
        RECT 6.4 0 6.65 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 3.5 4.4 3.8 ;
        RECT 1.5 3.5 2 3.8 ;
      LAYER MET2 ;
        RECT 3.9 3.45 4.4 3.85 ;
        RECT 1.5 3.5 4.4 3.8 ;
        RECT 1.5 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.62 3.52 1.88 3.78 ;
        RECT 4.02 3.52 4.28 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 2.85 5.7 3.15 ;
        RECT 2.35 2.85 2.85 3.15 ;
      LAYER MET2 ;
        RECT 5.2 2.8 5.7 3.2 ;
        RECT 2.35 2.85 5.7 3.15 ;
        RECT 2.35 2.8 2.85 3.2 ;
      LAYER VIA12 ;
        RECT 2.47 2.87 2.73 3.13 ;
        RECT 5.32 2.87 5.58 3.13 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
        RECT 0.55 0.95 0.8 7.15 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.2 4.8 7.7 5.1 ;
        RECT 7.25 4.75 7.6 5.15 ;
        RECT 7.25 0.95 7.5 7.15 ;
      LAYER MET2 ;
        RECT 7.2 4.75 7.7 5.15 ;
      LAYER VIA12 ;
        RECT 7.32 4.82 7.58 5.08 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 6.05 4.75 6.55 5.15 ;
      RECT 3 4.75 3.5 5.15 ;
      RECT 3 4.8 6.55 5.1 ;
    LAYER VIA12 ;
      RECT 6.17 4.82 6.43 5.08 ;
      RECT 3.12 4.82 3.38 5.08 ;
    LAYER MET1 ;
      RECT 5.55 3.5 5.8 7.15 ;
      RECT 5.55 3.5 7 3.8 ;
      RECT 4.7 3.5 7 3.75 ;
      RECT 4.7 1.35 4.95 3.75 ;
      RECT 5.55 0.85 5.8 1.9 ;
      RECT 3.85 0.85 4.1 1.9 ;
      RECT 3.85 0.85 5.8 1.1 ;
      RECT 2.25 4.8 2.5 7.15 ;
      RECT 1.05 4.8 3.5 5.1 ;
      RECT 3.1 0.95 3.35 5.1 ;
      RECT 6.05 4.8 6.55 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addh_1

MACRO gf180mcu_osu_sc_gp12t3v3__and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__and2_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.1 0 2.5 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 2.85 2.4 3.15 ;
      LAYER MET2 ;
        RECT 1.9 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.02 2.87 2.28 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 4.85 3.6 5.15 ;
        RECT 3.1 4.8 3.5 5.15 ;
        RECT 3.1 4.8 3.45 5.2 ;
        RECT 3.1 0.95 3.35 7.15 ;
      LAYER MET2 ;
        RECT 3.1 4.8 3.6 5.2 ;
      LAYER VIA12 ;
        RECT 3.22 4.87 3.48 5.13 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.35 4.1 2.85 4.5 ;
      RECT 1.3 4.1 1.8 4.5 ;
    LAYER VIA12 ;
      RECT 2.47 4.17 2.73 4.43 ;
      RECT 1.42 4.17 1.68 4.43 ;
    LAYER MET1 ;
      RECT 1.4 1.9 1.65 7.15 ;
      RECT 1.3 4.15 2.85 4.45 ;
      RECT 0.7 1.9 1.65 2.15 ;
      RECT 0.7 0.95 0.95 2.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__and2_1

MACRO gf180mcu_osu_sc_gp12t3v3__aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi21_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 1.4 6.2 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.95 0 3.2 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 4.15 2.1 4.45 ;
      LAYER MET2 ;
        RECT 1.6 4.1 2.1 4.5 ;
      LAYER VIA12 ;
        RECT 1.72 4.17 1.98 4.43 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 3.5 2.85 3.8 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.8 3.5 5.1 ;
        RECT 3.1 2.55 3.35 7.15 ;
        RECT 2.1 2.55 3.35 2.8 ;
        RECT 2.1 0.95 2.35 2.8 ;
      LAYER MET2 ;
        RECT 3 4.75 3.5 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 4.82 3.38 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.25 5.7 2.5 7.15 ;
      RECT 0.55 5.7 0.8 7.15 ;
      RECT 0.55 5.7 2.5 5.95 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi21_1

MACRO gf180mcu_osu_sc_gp12t3v3__aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi22_1 0 0 ;
  SIZE 5.35 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.35 8.1 ;
        RECT 1.4 6.2 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.35 0.6 ;
        RECT 3.5 0 3.75 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 4.15 2.1 4.45 ;
      LAYER MET2 ;
        RECT 1.6 4.1 2.1 4.5 ;
      LAYER VIA12 ;
        RECT 1.72 4.17 1.98 4.43 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 3.5 2.85 3.8 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 4.15 3.8 4.45 ;
      LAYER MET2 ;
        RECT 3.3 4.1 3.8 4.5 ;
      LAYER VIA12 ;
        RECT 3.42 4.17 3.68 4.43 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.3 4.8 4.8 5.1 ;
        RECT 4.45 6 4.75 6.5 ;
        RECT 4.45 4.8 4.7 6.5 ;
        RECT 4.4 3 4.65 5.1 ;
        RECT 2.1 3 4.65 3.25 ;
        RECT 2.1 0.95 2.35 3.25 ;
        RECT 3 6.1 3.5 6.4 ;
        RECT 3.1 6.1 3.35 7.15 ;
      LAYER MET2 ;
        RECT 4.35 6.05 4.85 6.45 ;
        RECT 3 6.1 4.85 6.4 ;
        RECT 3 6.05 3.5 6.45 ;
        RECT 4.3 4.75 4.8 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 6.12 3.38 6.38 ;
        RECT 4.42 4.82 4.68 5.08 ;
        RECT 4.47 6.12 4.73 6.38 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.95 5.6 4.2 7.15 ;
      RECT 2.25 5.6 2.5 7.15 ;
      RECT 0.55 5.6 0.8 7.15 ;
      RECT 0.55 5.6 4.2 5.85 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi22_1

MACRO gf180mcu_osu_sc_gp12t3v3__buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_1 0 0 ;
  SIZE 3.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.1 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.1 0.6 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 4.8 2.65 5.1 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.15 4.75 2.65 5.15 ;
      LAYER VIA12 ;
        RECT 2.27 4.82 2.53 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_1

MACRO gf180mcu_osu_sc_gp12t3v3__buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_16 0 0 ;
  SIZE 15.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15.8 8.1 ;
        RECT 15 5.45 15.25 8.1 ;
        RECT 13.3 5.45 13.55 8.1 ;
        RECT 11.6 5.45 11.85 8.1 ;
        RECT 9.9 5.45 10.15 8.1 ;
        RECT 8.2 5.45 8.45 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.05 4.8 14.55 5.1 ;
        RECT 14.15 0.95 14.4 7.15 ;
        RECT 2.25 4.85 14.4 5.15 ;
        RECT 2.25 2.05 14.4 2.3 ;
        RECT 12.45 0.95 12.7 7.15 ;
        RECT 10.75 0.95 11 7.15 ;
        RECT 9.05 0.95 9.3 7.15 ;
        RECT 7.35 0.95 7.6 7.15 ;
        RECT 5.65 0.95 5.9 7.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 14 4.85 14.55 5.15 ;
        RECT 14.05 4.75 14.55 5.15 ;
      LAYER VIA12 ;
        RECT 14.17 4.82 14.43 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_16

MACRO gf180mcu_osu_sc_gp12t3v3__buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_2 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 4.8 2.65 5.1 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.15 4.75 2.65 5.15 ;
      LAYER VIA12 ;
        RECT 2.27 4.82 2.53 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_2

MACRO gf180mcu_osu_sc_gp12t3v3__buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_4 0 0 ;
  SIZE 5.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.6 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.6 0.6 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.85 4.8 4.35 5.1 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 4.85 4.2 5.15 ;
        RECT 2.25 2.05 4.2 2.3 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 3.8 4.85 4.35 5.15 ;
        RECT 3.85 4.75 4.35 5.15 ;
      LAYER VIA12 ;
        RECT 3.97 4.82 4.23 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_4

MACRO gf180mcu_osu_sc_gp12t3v3__buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_8 0 0 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 9 8.1 ;
        RECT 8.2 5.45 8.45 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9 0.6 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 4.8 7.75 5.1 ;
        RECT 7.35 0.95 7.6 7.15 ;
        RECT 2.25 4.85 7.6 5.15 ;
        RECT 2.25 2.05 7.6 2.3 ;
        RECT 5.65 0.95 5.9 7.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 7.2 4.85 7.75 5.15 ;
        RECT 7.25 4.75 7.75 5.15 ;
      LAYER VIA12 ;
        RECT 7.37 4.82 7.63 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_8

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_1 0 0 ;
  SIZE 3.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.1 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.1 0.6 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 4.8 2.65 5.1 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.15 4.75 2.65 5.15 ;
      LAYER VIA12 ;
        RECT 2.27 4.82 2.53 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_1

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_16 0 0 ;
  SIZE 15.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15.8 8.1 ;
        RECT 15 5.45 15.25 8.1 ;
        RECT 13.3 5.45 13.55 8.1 ;
        RECT 11.6 5.45 11.85 8.1 ;
        RECT 9.9 5.45 10.15 8.1 ;
        RECT 8.2 5.45 8.45 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 4.85 14.55 5.15 ;
        RECT 14.15 0.95 14.4 7.15 ;
        RECT 2.25 2.05 14.4 2.3 ;
        RECT 12.45 0.95 12.7 7.15 ;
        RECT 10.75 0.95 11 7.15 ;
        RECT 9.05 0.95 9.3 7.15 ;
        RECT 7.35 0.95 7.6 7.15 ;
        RECT 5.65 0.95 5.9 7.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 14.05 4.8 14.55 5.2 ;
        RECT 14 4.85 14.55 5.15 ;
      LAYER VIA12 ;
        RECT 14.17 4.87 14.43 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_16

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_2 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 4.85 2.65 5.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.15 4.8 2.65 5.2 ;
      LAYER VIA12 ;
        RECT 2.27 4.87 2.53 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_2

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_4 0 0 ;
  SIZE 5.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.6 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.6 0.6 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 4.85 4.35 5.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 2.05 4.2 2.3 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 3.85 4.8 4.35 5.2 ;
        RECT 3.8 4.85 4.35 5.15 ;
      LAYER VIA12 ;
        RECT 3.97 4.87 4.23 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_4

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_8 0 0 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 9 8.1 ;
        RECT 8.2 5.45 8.45 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9 0.6 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 4.85 7.75 5.15 ;
        RECT 7.35 0.95 7.6 7.15 ;
        RECT 2.25 2.05 7.6 2.3 ;
        RECT 5.65 0.95 5.9 7.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 7.25 4.8 7.75 5.2 ;
        RECT 7.2 4.85 7.75 5.15 ;
      LAYER VIA12 ;
        RECT 7.37 4.87 7.63 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_8

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_1 0 0 ;
  SIZE 2.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.2 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_1

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_16 0 0 ;
  SIZE 15 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15 8.1 ;
        RECT 14.15 5.45 14.4 8.1 ;
        RECT 12.45 5.45 12.7 8.1 ;
        RECT 10.75 5.45 11 8.1 ;
        RECT 9.05 5.45 9.3 8.1 ;
        RECT 7.35 5.45 7.6 8.1 ;
        RECT 5.65 5.45 5.9 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15 0.6 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 12.45 0 12.7 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 9.05 0 9.3 1.8 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.3 0.95 13.55 7.15 ;
        RECT 1.4 4.45 13.55 4.7 ;
        RECT 13.15 4.35 13.55 4.7 ;
        RECT 1.4 2.05 13.55 2.3 ;
        RECT 11.6 0.95 11.85 7.15 ;
        RECT 9.9 0.95 10.15 7.15 ;
        RECT 8.2 0.95 8.45 7.15 ;
        RECT 6.5 0.95 6.75 7.15 ;
        RECT 4.8 0.95 5.05 7.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 13.15 4.35 13.65 4.75 ;
      LAYER VIA12 ;
        RECT 13.27 4.42 13.53 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_16

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_2 0 0 ;
  SIZE 3.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.2 8.1 ;
        RECT 2.3 5.45 2.55 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 3.5 1.15 3.8 ;
      LAYER MET2 ;
        RECT 0.65 3.45 1.15 3.85 ;
      LAYER VIA12 ;
        RECT 0.77 3.52 1.03 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 4.4 2 4.7 ;
        RECT 1.4 4.25 1.85 4.8 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 1.5 4.35 2 4.75 ;
      LAYER VIA12 ;
        RECT 1.62 4.42 1.88 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_2

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_4 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 4.45 3.35 4.7 ;
        RECT 2.95 4.35 3.35 4.7 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 2.95 4.35 3.45 4.75 ;
      LAYER VIA12 ;
        RECT 3.07 4.42 3.33 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_4

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_8 0 0 ;
  SIZE 8.15 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 8.15 8.1 ;
        RECT 7.35 5.45 7.6 8.1 ;
        RECT 5.65 5.45 5.9 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.15 0.6 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.5 0.95 6.75 7.15 ;
        RECT 1.4 4.45 6.75 4.7 ;
        RECT 6.35 4.35 6.75 4.7 ;
        RECT 1.4 2.05 6.75 2.3 ;
        RECT 4.8 0.95 5.05 7.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 6.35 4.35 6.85 4.75 ;
      LAYER VIA12 ;
        RECT 6.47 4.42 6.73 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_8

MACRO gf180mcu_osu_sc_gp12t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dff_1 0 0 ;
  SIZE 13 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 13 8.1 ;
        RECT 11.3 5.45 11.55 8.1 ;
        RECT 8.85 5.45 9.1 8.1 ;
        RECT 7.25 6.2 7.5 8.1 ;
        RECT 4.45 5.45 4.7 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 13 0.6 ;
        RECT 11.3 0 11.55 1.8 ;
        RECT 8.85 0 9.1 1.45 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 4.45 0 4.7 1.4 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.65 4.15 8.15 4.45 ;
        RECT 5.5 4.15 6.55 4.45 ;
        RECT 5.4 2.15 5.9 2.45 ;
        RECT 5.5 2.15 5.8 4.45 ;
        RECT 2.6 4.15 3.75 4.45 ;
        RECT 3.25 2.2 3.75 2.5 ;
        RECT 3.35 2.2 3.65 4.45 ;
      LAYER MET2 ;
        RECT 3.25 4.15 8.15 4.45 ;
        RECT 7.7 4.1 8.1 4.5 ;
        RECT 6.05 4.1 6.55 4.5 ;
        RECT 3.25 4.1 3.7 4.5 ;
      LAYER VIA12 ;
        RECT 3.37 4.17 3.63 4.43 ;
        RECT 6.17 4.17 6.43 4.43 ;
        RECT 7.77 4.17 8.03 4.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.5 2.4 3.8 ;
      LAYER MET2 ;
        RECT 1.75 3.5 2.55 3.8 ;
        RECT 1.9 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.02 3.52 2.28 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.15 4.8 12.65 5.15 ;
        RECT 12.15 4.75 12.6 5.15 ;
        RECT 12.15 0.95 12.4 7.15 ;
      LAYER MET2 ;
        RECT 12.15 4.8 12.65 5.1 ;
        RECT 12.2 4.75 12.6 5.15 ;
      LAYER VIA12 ;
        RECT 12.27 4.82 12.53 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.45 4.15 11.9 4.45 ;
        RECT 11.55 2.05 11.8 4.45 ;
        RECT 10.45 2.05 11.8 2.3 ;
        RECT 10.45 4.15 10.7 7.15 ;
        RECT 10.45 0.95 10.7 2.3 ;
      LAYER MET2 ;
        RECT 11.4 4.15 11.9 4.45 ;
        RECT 11.45 4.1 11.85 4.5 ;
      LAYER VIA12 ;
        RECT 11.52 4.17 11.78 4.43 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 6.75 4.75 7.15 5.15 ;
      RECT 6.7 4.8 9.9 5.1 ;
      RECT 9.6 2.85 9.9 5.1 ;
      RECT 10.7 2.8 11.1 3.2 ;
      RECT 9.6 2.85 11.15 3.15 ;
      RECT 9 1.65 9.4 2.05 ;
      RECT 8.5 1.7 9.45 2 ;
      RECT 5.8 1.5 6.2 1.9 ;
      RECT 5.75 1.55 8.8 1.85 ;
      RECT 5.75 1.65 9.4 1.85 ;
      RECT 8.05 2.8 8.45 3.2 ;
      RECT 6.1 2.8 6.5 3.2 ;
      RECT 6.05 2.85 8.55 3.15 ;
      RECT 6.8 3.45 7.2 3.85 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.1 2.15 4.5 2.55 ;
      RECT 0.45 2.15 0.85 2.55 ;
      RECT 0.4 2.2 4.55 2.5 ;
    LAYER VIA12 ;
      RECT 10.77 2.87 11.03 3.13 ;
      RECT 9.07 1.72 9.33 1.98 ;
      RECT 8.12 2.87 8.38 3.13 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.82 4.82 7.08 5.08 ;
      RECT 6.17 2.87 6.43 3.13 ;
      RECT 5.87 1.57 6.13 1.83 ;
      RECT 4.17 2.22 4.43 2.48 ;
      RECT 0.52 2.22 0.78 2.48 ;
    LAYER MET1 ;
      RECT 9.7 0.95 9.95 7.15 ;
      RECT 9.7 2.85 11.15 3.15 ;
      RECT 9.05 1.7 9.35 3.25 ;
      RECT 8.95 2.85 9.45 3.15 ;
      RECT 8.95 1.7 9.45 2 ;
      RECT 8.1 4.75 8.35 7.15 ;
      RECT 8.1 4.75 8.9 5 ;
      RECT 8.6 3.55 8.9 5 ;
      RECT 8.1 3.55 8.9 3.8 ;
      RECT 8.1 2.75 8.4 3.8 ;
      RECT 8.1 0.95 8.35 3.8 ;
      RECT 6.7 4.8 7.2 5.1 ;
      RECT 6.8 3.45 7.1 5.1 ;
      RECT 6.75 3.5 7.3 3.8 ;
      RECT 6.8 3.45 7.2 3.8 ;
      RECT 5.85 5.95 6.1 7.15 ;
      RECT 4.95 5.95 6.1 6.2 ;
      RECT 4.95 3.45 5.2 6.2 ;
      RECT 4.9 1.6 5.15 3.7 ;
      RECT 4.9 1.6 6.25 1.85 ;
      RECT 5.85 1.55 6.25 1.85 ;
      RECT 5.85 0.95 6.1 1.85 ;
      RECT 4.05 4.8 4.55 5.1 ;
      RECT 4.15 2.2 4.45 5.1 ;
      RECT 4.05 2.2 4.55 2.5 ;
      RECT 3.05 4.95 3.3 7.15 ;
      RECT 1.4 4.95 3.3 5.2 ;
      RECT 1.4 2.25 1.65 5.2 ;
      RECT 1.05 4.15 1.65 4.45 ;
      RECT 1.4 2.25 2.4 2.5 ;
      RECT 2 1.55 2.4 2.5 ;
      RECT 2 1.55 3.3 1.8 ;
      RECT 3.05 0.95 3.3 1.8 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.5 2.1 0.8 2.6 ;
      RECT 6.05 2.85 6.55 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dff_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffn_1 0 0 ;
  SIZE 14.25 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 14.25 8.1 ;
        RECT 12.55 5.45 12.8 8.1 ;
        RECT 9.95 5.45 10.35 8.1 ;
        RECT 7.25 6.2 7.5 8.1 ;
        RECT 4.45 5.45 4.7 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.25 0.6 ;
        RECT 12.55 0 12.8 1.8 ;
        RECT 9.95 0 10.35 1.45 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 4.45 0 4.7 1.4 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9.5 2.85 10 3.15 ;
        RECT 9.6 2.75 9.9 3.25 ;
      LAYER MET2 ;
        RECT 9.5 2.85 10 3.15 ;
        RECT 9.55 2.8 9.95 3.2 ;
      LAYER VIA12 ;
        RECT 9.62 2.87 9.88 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.5 2.4 3.8 ;
      LAYER MET2 ;
        RECT 1.75 3.5 2.55 3.8 ;
        RECT 1.9 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.02 3.52 2.28 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.4 4.8 13.9 5.15 ;
        RECT 13.4 4.75 13.85 5.15 ;
        RECT 13.4 0.95 13.65 7.15 ;
      LAYER MET2 ;
        RECT 13.4 4.8 13.9 5.1 ;
        RECT 13.45 4.75 13.85 5.15 ;
      LAYER VIA12 ;
        RECT 13.52 4.82 13.78 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.7 4.15 13.15 4.45 ;
        RECT 12.8 2.05 13.05 4.45 ;
        RECT 11.7 2.05 13.05 2.3 ;
        RECT 11.7 4.15 11.95 7.15 ;
        RECT 11.7 0.95 11.95 2.3 ;
      LAYER MET2 ;
        RECT 12.65 4.15 13.15 4.45 ;
        RECT 12.7 4.1 13.1 4.5 ;
      LAYER VIA12 ;
        RECT 12.77 4.17 13.03 4.43 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 6.75 4.75 7.15 5.15 ;
      RECT 6.7 4.8 11.15 5.1 ;
      RECT 10.85 2.85 11.15 5.1 ;
      RECT 11.95 2.8 12.35 3.2 ;
      RECT 10.85 2.85 12.4 3.15 ;
      RECT 10.25 1.65 10.65 2.05 ;
      RECT 9.5 1.7 10.7 2 ;
      RECT 5.8 1.5 6.2 1.9 ;
      RECT 5.75 1.55 9.9 1.85 ;
      RECT 5.75 1.65 10.65 1.85 ;
      RECT 8.9 4.1 9.3 4.5 ;
      RECT 7.7 4.1 8.1 4.5 ;
      RECT 6.05 4.1 6.55 4.5 ;
      RECT 3.25 4.1 3.7 4.5 ;
      RECT 3.25 4.15 9.35 4.45 ;
      RECT 8.05 2.8 8.45 3.2 ;
      RECT 6.1 2.8 6.5 3.2 ;
      RECT 6.05 2.85 8.55 3.15 ;
      RECT 6.8 3.45 7.2 3.85 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.1 2.15 4.5 2.55 ;
      RECT 0.45 2.15 0.85 2.55 ;
      RECT 0.4 2.2 4.55 2.5 ;
    LAYER VIA12 ;
      RECT 12.02 2.87 12.28 3.13 ;
      RECT 10.32 1.72 10.58 1.98 ;
      RECT 8.97 4.17 9.23 4.43 ;
      RECT 8.12 2.87 8.38 3.13 ;
      RECT 7.77 4.17 8.03 4.43 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.82 4.82 7.08 5.08 ;
      RECT 6.17 2.87 6.43 3.13 ;
      RECT 6.17 4.17 6.43 4.43 ;
      RECT 5.87 1.57 6.13 1.83 ;
      RECT 4.17 2.22 4.43 2.48 ;
      RECT 3.37 4.17 3.63 4.43 ;
      RECT 0.52 2.22 0.78 2.48 ;
    LAYER MET1 ;
      RECT 10.95 0.95 11.2 7.15 ;
      RECT 10.95 2.85 12.4 3.15 ;
      RECT 10.3 1.7 10.6 5.2 ;
      RECT 10.2 4.8 10.7 5.1 ;
      RECT 10.2 1.7 10.7 2 ;
      RECT 9.1 5.45 9.35 7.15 ;
      RECT 8.95 1.6 9.25 5.7 ;
      RECT 9.1 0.95 9.35 1.85 ;
      RECT 8.1 4.75 8.35 7.15 ;
      RECT 8.1 4.75 8.7 5 ;
      RECT 8.4 3.55 8.7 5 ;
      RECT 8.1 2.75 8.4 3.8 ;
      RECT 8.1 0.95 8.35 3.8 ;
      RECT 6.7 4.8 7.2 5.1 ;
      RECT 6.8 3.5 7.1 5.1 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 5.5 4.15 6.55 4.45 ;
      RECT 5.5 2.15 5.8 4.45 ;
      RECT 5.4 2.15 5.9 2.45 ;
      RECT 5.85 5.95 6.1 7.15 ;
      RECT 4.95 5.95 6.1 6.2 ;
      RECT 4.95 3.45 5.2 6.2 ;
      RECT 4.9 1.6 5.15 3.7 ;
      RECT 4.9 1.6 6.25 1.85 ;
      RECT 5.85 1.55 6.25 1.85 ;
      RECT 5.85 0.95 6.1 1.85 ;
      RECT 4.05 4.8 4.55 5.1 ;
      RECT 4.15 2.2 4.45 5.1 ;
      RECT 4.05 2.2 4.55 2.5 ;
      RECT 2.6 4.15 3.75 4.45 ;
      RECT 3.35 2.2 3.65 4.45 ;
      RECT 3.25 2.2 3.75 2.5 ;
      RECT 3.05 4.95 3.3 7.15 ;
      RECT 1.4 4.95 3.3 5.2 ;
      RECT 1.4 2.25 1.65 5.2 ;
      RECT 1.05 4.15 1.65 4.45 ;
      RECT 1.4 2.25 2.4 2.5 ;
      RECT 2 1.55 2.4 2.5 ;
      RECT 2 1.55 3.3 1.8 ;
      RECT 3.05 0.95 3.3 1.8 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.5 2.1 0.8 2.6 ;
      RECT 7.65 4.15 8.15 4.45 ;
      RECT 6.05 2.85 6.55 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffr_1 0 0 ;
  SIZE 17.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 17.6 8.1 ;
        RECT 15.95 5.45 16.2 8.1 ;
        RECT 12.95 5.45 13.2 8.1 ;
        RECT 10.75 6.2 11 8.1 ;
        RECT 7.95 5.45 8.2 8.1 ;
        RECT 4.9 5.45 5.15 8.1 ;
        RECT 3.55 5.45 3.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 17.6 0.6 ;
        RECT 15.95 0 16.2 1.8 ;
        RECT 14.2 0 14.45 1.8 ;
        RECT 12.5 0 12.75 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 7.95 0 8.2 1.4 ;
        RECT 4.9 0 5.15 1.8 ;
        RECT 4 0 4.25 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 11.15 4.15 11.65 4.45 ;
        RECT 9 4.15 10.05 4.45 ;
        RECT 8.9 2.15 9.4 2.45 ;
        RECT 9 2.15 9.3 4.45 ;
        RECT 6.1 4.15 7.25 4.45 ;
        RECT 6.75 2.2 7.25 2.5 ;
        RECT 6.85 2.2 7.15 4.45 ;
      LAYER MET2 ;
        RECT 6.75 4.15 11.65 4.45 ;
        RECT 11.2 4.1 11.6 4.5 ;
        RECT 9.55 4.1 10.05 4.5 ;
        RECT 6.75 4.1 7.2 4.5 ;
      LAYER VIA12 ;
        RECT 6.87 4.17 7.13 4.43 ;
        RECT 9.67 4.17 9.93 4.43 ;
        RECT 11.27 4.17 11.53 4.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.4 3.5 5.9 3.8 ;
      LAYER MET2 ;
        RECT 5.4 3.45 5.9 3.85 ;
      LAYER VIA12 ;
        RECT 5.52 3.52 5.78 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.8 4.8 17.3 5.15 ;
        RECT 16.8 4.75 17.25 5.15 ;
        RECT 16.8 0.95 17.05 7.15 ;
      LAYER MET2 ;
        RECT 16.8 4.8 17.3 5.1 ;
        RECT 16.85 4.75 17.25 5.15 ;
      LAYER VIA12 ;
        RECT 16.92 4.82 17.18 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.1 4.15 16.55 4.45 ;
        RECT 16.2 2.05 16.45 4.45 ;
        RECT 15.1 2.05 16.45 2.3 ;
        RECT 15.1 4.15 15.35 7.15 ;
        RECT 15.1 0.95 15.35 2.3 ;
      LAYER MET2 ;
        RECT 16.05 4.15 16.55 4.45 ;
        RECT 16.1 4.1 16.5 4.5 ;
      LAYER VIA12 ;
        RECT 16.17 4.17 16.43 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  OBS
    LAYER MET2 ;
      RECT 15.35 2.8 15.75 3.2 ;
      RECT 15 2.85 15.8 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 13.75 2.1 14.35 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 13.75 0.9 14.05 2.5 ;
      RECT 2.75 0.9 14.05 1.2 ;
      RECT 12.4 2.1 12.9 2.5 ;
      RECT 12.4 1.55 12.8 2.5 ;
      RECT 9.3 1.5 9.7 1.9 ;
      RECT 9.25 1.55 12.8 1.85 ;
      RECT 12.45 4.75 12.85 5.15 ;
      RECT 10.25 4.75 10.65 5.15 ;
      RECT 10.2 4.8 12.9 5.1 ;
      RECT 11.55 2.8 11.95 3.2 ;
      RECT 9.6 2.8 10 3.2 ;
      RECT 9.55 2.85 12.05 3.15 ;
      RECT 10.3 3.45 10.7 3.85 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 7.6 2.15 8 2.55 ;
      RECT 3.85 2.15 4.35 2.55 ;
      RECT 3.85 2.2 8.05 2.5 ;
      RECT 14.25 4.75 14.75 5.15 ;
    LAYER VIA12 ;
      RECT 15.42 2.87 15.68 3.13 ;
      RECT 14.37 4.82 14.63 5.08 ;
      RECT 13.97 2.17 14.23 2.43 ;
      RECT 12.52 2.17 12.78 2.43 ;
      RECT 12.52 4.82 12.78 5.08 ;
      RECT 11.62 2.87 11.88 3.13 ;
      RECT 10.37 3.52 10.63 3.78 ;
      RECT 10.32 4.82 10.58 5.08 ;
      RECT 9.67 2.87 9.93 3.13 ;
      RECT 9.37 1.57 9.63 1.83 ;
      RECT 7.67 2.22 7.93 2.48 ;
      RECT 3.97 2.22 4.23 2.48 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 14.35 2.85 14.6 7.15 ;
      RECT 12.5 4.7 12.8 5.2 ;
      RECT 12.5 4.8 14.75 5.1 ;
      RECT 13.35 2.85 15.8 3.15 ;
      RECT 13.35 0.95 13.6 3.15 ;
      RECT 11.6 4.75 11.85 7.15 ;
      RECT 11.6 4.75 12.15 5 ;
      RECT 11.9 3.55 12.15 5 ;
      RECT 11.6 2.75 11.9 3.8 ;
      RECT 11.6 0.95 11.85 3.8 ;
      RECT 10.2 4.8 10.7 5.1 ;
      RECT 10.3 3.5 10.6 5.1 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 9.35 5.95 9.6 7.15 ;
      RECT 8.45 5.95 9.6 6.2 ;
      RECT 8.45 3.45 8.7 6.2 ;
      RECT 8.4 1.6 8.65 3.7 ;
      RECT 8.4 1.6 9.75 1.85 ;
      RECT 9.35 1.55 9.75 1.85 ;
      RECT 9.35 0.95 9.6 1.85 ;
      RECT 7.55 4.8 8.05 5.1 ;
      RECT 7.65 2.2 7.95 5.1 ;
      RECT 7.55 2.2 8.05 2.5 ;
      RECT 6.55 4.95 6.8 7.15 ;
      RECT 4.9 4.95 6.8 5.2 ;
      RECT 4.9 2.25 5.15 5.2 ;
      RECT 3.85 4.15 5.15 4.45 ;
      RECT 4.9 2.25 5.9 2.5 ;
      RECT 5.5 1.55 5.9 2.5 ;
      RECT 5.5 1.55 6.8 1.8 ;
      RECT 6.55 0.95 6.8 1.8 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 3.95 2.15 4.2 2.55 ;
      RECT 3 2.2 4.35 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 13.85 2.15 14.35 2.45 ;
      RECT 12.4 2.15 12.9 2.45 ;
      RECT 9.55 2.85 10.05 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffr_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffrn_1 0 0 ;
  SIZE 19.25 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 19.25 8.1 ;
        RECT 17.6 5.45 17.85 8.1 ;
        RECT 14.6 5.45 14.85 8.1 ;
        RECT 13.4 5.45 13.65 8.1 ;
        RECT 10.75 6.2 11 8.1 ;
        RECT 7.95 5.45 8.2 8.1 ;
        RECT 4.9 5.45 5.15 8.1 ;
        RECT 3.55 5.45 3.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 19.25 0.6 ;
        RECT 17.6 0 17.85 1.8 ;
        RECT 15.85 0 16.1 1.8 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 13.4 0 13.65 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 7.95 0 8.2 1.4 ;
        RECT 4.9 0 5.15 1.8 ;
        RECT 4 0 4.25 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 13.15 2.85 13.65 3.15 ;
      LAYER MET2 ;
        RECT 13.15 2.8 13.65 3.2 ;
      LAYER VIA12 ;
        RECT 13.27 2.87 13.53 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.4 3.5 5.9 3.8 ;
      LAYER MET2 ;
        RECT 5.4 3.45 5.9 3.85 ;
      LAYER VIA12 ;
        RECT 5.52 3.52 5.78 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 18.45 4.8 18.95 5.15 ;
        RECT 18.45 4.75 18.9 5.15 ;
        RECT 18.45 0.95 18.7 7.15 ;
      LAYER MET2 ;
        RECT 18.45 4.8 18.95 5.1 ;
        RECT 18.5 4.75 18.9 5.15 ;
      LAYER VIA12 ;
        RECT 18.57 4.82 18.83 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.75 4.15 18.2 4.45 ;
        RECT 17.85 2.05 18.1 4.45 ;
        RECT 16.75 2.05 18.1 2.3 ;
        RECT 16.75 4.15 17 7.15 ;
        RECT 16.75 0.95 17 2.3 ;
      LAYER MET2 ;
        RECT 17.7 4.15 18.2 4.45 ;
        RECT 17.75 4.1 18.15 4.5 ;
      LAYER VIA12 ;
        RECT 17.82 4.17 18.08 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  OBS
    LAYER MET2 ;
      RECT 17 2.8 17.4 3.2 ;
      RECT 16.65 2.85 17.45 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 15.4 2.1 16 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 15.4 0.9 15.7 2.5 ;
      RECT 2.75 0.9 15.7 1.2 ;
      RECT 14.05 2.1 14.55 2.5 ;
      RECT 14.05 1.55 14.45 2.5 ;
      RECT 9.3 1.5 9.7 1.9 ;
      RECT 9.25 1.55 14.45 1.85 ;
      RECT 14.1 4.75 14.5 5.15 ;
      RECT 10.25 4.75 10.65 5.15 ;
      RECT 10.2 4.8 14.55 5.1 ;
      RECT 12.45 4.1 12.9 4.5 ;
      RECT 11.2 4.1 11.6 4.5 ;
      RECT 9.55 4.1 10.05 4.5 ;
      RECT 6.75 4.1 7.2 4.5 ;
      RECT 6.75 4.15 12.9 4.45 ;
      RECT 11.55 2.8 11.95 3.2 ;
      RECT 9.6 2.8 10 3.2 ;
      RECT 9.55 2.85 12.05 3.15 ;
      RECT 10.3 3.45 10.7 3.85 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 7.6 2.15 8 2.55 ;
      RECT 3.85 2.15 4.35 2.55 ;
      RECT 3.85 2.2 8.05 2.5 ;
      RECT 15.9 4.75 16.4 5.15 ;
    LAYER VIA12 ;
      RECT 17.07 2.87 17.33 3.13 ;
      RECT 16.02 4.82 16.28 5.08 ;
      RECT 15.62 2.17 15.88 2.43 ;
      RECT 14.17 2.17 14.43 2.43 ;
      RECT 14.17 4.82 14.43 5.08 ;
      RECT 12.52 4.17 12.78 4.43 ;
      RECT 11.62 2.87 11.88 3.13 ;
      RECT 11.27 4.17 11.53 4.43 ;
      RECT 10.37 3.52 10.63 3.78 ;
      RECT 10.32 4.82 10.58 5.08 ;
      RECT 9.67 2.87 9.93 3.13 ;
      RECT 9.67 4.17 9.93 4.43 ;
      RECT 9.37 1.57 9.63 1.83 ;
      RECT 7.67 2.22 7.93 2.48 ;
      RECT 6.87 4.17 7.13 4.43 ;
      RECT 3.97 2.22 4.23 2.48 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 16 2.85 16.25 7.15 ;
      RECT 14.15 4.7 14.45 5.2 ;
      RECT 14.15 4.8 16.4 5.1 ;
      RECT 15 2.85 17.45 3.15 ;
      RECT 15 0.95 15.25 3.15 ;
      RECT 12.55 0.95 12.8 7.15 ;
      RECT 12.4 4.15 12.9 4.45 ;
      RECT 11.6 4.75 11.85 7.15 ;
      RECT 11.6 4.75 12.15 5 ;
      RECT 11.9 3.55 12.15 5 ;
      RECT 11.6 2.75 11.9 3.8 ;
      RECT 11.6 0.95 11.85 3.8 ;
      RECT 10.2 4.8 10.7 5.1 ;
      RECT 10.3 3.5 10.6 5.1 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 9 4.15 10.05 4.45 ;
      RECT 9 2.15 9.3 4.45 ;
      RECT 8.9 2.15 9.4 2.45 ;
      RECT 9.35 5.95 9.6 7.15 ;
      RECT 8.45 5.95 9.6 6.2 ;
      RECT 8.45 3.45 8.7 6.2 ;
      RECT 8.4 1.6 8.65 3.7 ;
      RECT 8.4 1.6 9.75 1.85 ;
      RECT 9.35 1.55 9.75 1.85 ;
      RECT 9.35 0.95 9.6 1.85 ;
      RECT 7.55 4.8 8.05 5.1 ;
      RECT 7.65 2.2 7.95 5.1 ;
      RECT 7.55 2.2 8.05 2.5 ;
      RECT 6.1 4.15 7.25 4.45 ;
      RECT 6.85 2.2 7.15 4.45 ;
      RECT 6.75 2.2 7.25 2.5 ;
      RECT 6.55 4.95 6.8 7.15 ;
      RECT 4.9 4.95 6.8 5.2 ;
      RECT 4.9 2.25 5.15 5.2 ;
      RECT 3.85 4.15 5.15 4.45 ;
      RECT 4.9 2.25 5.9 2.5 ;
      RECT 5.5 1.55 5.9 2.5 ;
      RECT 5.5 1.55 6.8 1.8 ;
      RECT 6.55 0.95 6.8 1.8 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 3.95 2.15 4.2 2.55 ;
      RECT 3 2.2 4.35 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 15.5 2.15 16 2.45 ;
      RECT 14.05 2.15 14.55 2.45 ;
      RECT 11.15 4.15 11.65 4.45 ;
      RECT 9.55 2.85 10.05 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffrn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffs_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffs_1 0 0 ;
  SIZE 15.45 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15.45 8.1 ;
        RECT 13.8 5.45 14.05 8.1 ;
        RECT 11.35 6.7 11.6 8.1 ;
        RECT 8.9 6.2 9.15 8.1 ;
        RECT 6.1 5.45 6.35 8.1 ;
        RECT 3.05 5.45 3.3 8.1 ;
        RECT 1.45 6.2 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.45 0.6 ;
        RECT 13.8 0 14.05 1.8 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.9 0 9.15 1.8 ;
        RECT 6.1 0 6.35 1.4 ;
        RECT 3.05 0 3.3 1.8 ;
        RECT 2.15 0 2.4 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9.3 4.15 9.8 4.45 ;
        RECT 7.15 4.15 8.2 4.45 ;
        RECT 7.05 2.15 7.55 2.45 ;
        RECT 7.15 2.15 7.45 4.45 ;
        RECT 4.25 4.15 5.4 4.45 ;
        RECT 4.9 2.2 5.4 2.5 ;
        RECT 5 2.2 5.3 4.45 ;
      LAYER MET2 ;
        RECT 4.9 4.15 9.8 4.45 ;
        RECT 9.35 4.1 9.75 4.5 ;
        RECT 7.7 4.1 8.2 4.5 ;
        RECT 4.9 4.1 5.35 4.5 ;
      LAYER VIA12 ;
        RECT 5.02 4.17 5.28 4.43 ;
        RECT 7.82 4.17 8.08 4.43 ;
        RECT 9.42 4.17 9.68 4.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.55 3.5 4.05 3.8 ;
      LAYER MET2 ;
        RECT 3.55 3.45 4.05 3.85 ;
      LAYER VIA12 ;
        RECT 3.67 3.52 3.93 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.65 4.8 15.15 5.15 ;
        RECT 14.65 4.75 15.1 5.15 ;
        RECT 14.65 0.95 14.9 7.15 ;
      LAYER MET2 ;
        RECT 14.65 4.8 15.15 5.1 ;
        RECT 14.7 4.75 15.1 5.15 ;
      LAYER VIA12 ;
        RECT 14.77 4.82 15.03 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.95 4.15 14.4 4.45 ;
        RECT 14.05 2.05 14.3 4.45 ;
        RECT 12.95 2.05 14.3 2.3 ;
        RECT 12.95 4.15 13.2 7.15 ;
        RECT 12.95 0.95 13.2 2.3 ;
      LAYER MET2 ;
        RECT 13.9 4.15 14.4 4.45 ;
        RECT 13.95 4.1 14.35 4.5 ;
      LAYER VIA12 ;
        RECT 14.02 4.17 14.28 4.43 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.55 4.15 12.05 4.45 ;
        RECT 5.7 4.8 6.2 5.1 ;
        RECT 5.7 2.2 6.2 2.5 ;
        RECT 5.8 2.2 6.1 5.1 ;
        RECT 2.3 5.7 2.55 7.15 ;
        RECT 0.75 2.2 2.5 2.5 ;
        RECT 2.1 2.15 2.35 2.55 ;
        RECT 0.6 5.7 2.55 5.95 ;
        RECT 0.75 4.15 1.5 4.45 ;
        RECT 0.75 0.95 1 5.95 ;
        RECT 0.6 5.7 0.85 7.15 ;
      LAYER MET2 ;
        RECT 11.55 4.1 12.05 4.5 ;
        RECT 1.1 5.45 11.95 5.75 ;
        RECT 11.65 4.1 11.95 5.75 ;
        RECT 1 4.1 1.5 4.5 ;
        RECT 1.1 4.1 1.4 5.75 ;
        RECT 2 2.2 6.2 2.5 ;
        RECT 5.75 2.15 6.15 2.55 ;
        RECT 2 2.15 2.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.12 4.17 1.38 4.43 ;
        RECT 2.12 2.22 2.38 2.48 ;
        RECT 5.82 2.22 6.08 2.48 ;
        RECT 11.67 4.17 11.93 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 13.2 2.8 13.6 3.2 ;
      RECT 12.85 2.85 13.65 3.15 ;
      RECT 10.55 2.1 11.05 2.5 ;
      RECT 10.55 1.55 10.95 2.5 ;
      RECT 7.45 1.5 7.85 1.9 ;
      RECT 7.4 1.55 10.95 1.85 ;
      RECT 10.6 4.75 11 5.15 ;
      RECT 8.4 4.75 8.8 5.15 ;
      RECT 8.35 4.8 11.05 5.1 ;
      RECT 9.7 2.8 10.1 3.2 ;
      RECT 7.75 2.8 8.15 3.2 ;
      RECT 7.7 2.85 10.2 3.15 ;
      RECT 8.45 3.45 8.85 3.85 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 12.25 4.75 12.75 5.15 ;
      RECT 2 3.45 2.5 3.85 ;
    LAYER VIA12 ;
      RECT 13.27 2.87 13.53 3.13 ;
      RECT 12.37 4.82 12.63 5.08 ;
      RECT 10.67 2.17 10.93 2.43 ;
      RECT 10.67 4.82 10.93 5.08 ;
      RECT 9.77 2.87 10.03 3.13 ;
      RECT 8.52 3.52 8.78 3.78 ;
      RECT 8.47 4.82 8.73 5.08 ;
      RECT 7.82 2.87 8.08 3.13 ;
      RECT 7.52 1.57 7.78 1.83 ;
      RECT 2.12 3.52 2.38 3.78 ;
    LAYER MET1 ;
      RECT 12.35 2.85 12.65 5.2 ;
      RECT 10.65 4.7 10.95 5.2 ;
      RECT 10.65 4.8 12.65 5.1 ;
      RECT 12.05 2.85 13.65 3.15 ;
      RECT 12.05 0.95 12.3 3.15 ;
      RECT 12.2 6.2 12.45 7.15 ;
      RECT 10.5 6.2 10.75 7.15 ;
      RECT 10.5 6.2 12.45 6.45 ;
      RECT 9.75 4.75 10 7.15 ;
      RECT 9.75 4.75 10.3 5 ;
      RECT 10.05 3.55 10.3 5 ;
      RECT 9.75 2.75 10.05 3.8 ;
      RECT 9.75 0.95 10 3.8 ;
      RECT 8.35 4.8 8.85 5.1 ;
      RECT 8.45 3.5 8.75 5.1 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 7.5 5.95 7.75 7.15 ;
      RECT 6.6 5.95 7.75 6.2 ;
      RECT 6.6 3.45 6.85 6.2 ;
      RECT 6.55 1.6 6.8 3.7 ;
      RECT 6.55 1.6 7.9 1.85 ;
      RECT 7.5 1.55 7.9 1.85 ;
      RECT 7.5 0.95 7.75 1.85 ;
      RECT 4.7 4.95 4.95 7.15 ;
      RECT 3.05 4.95 4.95 5.2 ;
      RECT 3.05 2.25 3.3 5.2 ;
      RECT 2 3.5 3.3 3.8 ;
      RECT 3.05 2.25 4.05 2.5 ;
      RECT 3.65 1.55 4.05 2.5 ;
      RECT 3.65 1.55 4.95 1.8 ;
      RECT 4.7 0.95 4.95 1.8 ;
      RECT 10.55 2.15 11.05 2.45 ;
      RECT 7.7 2.85 8.2 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffs_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsn_1 0 0 ;
  SIZE 17.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 17.2 8.1 ;
        RECT 15.5 5.45 15.75 8.1 ;
        RECT 13.05 6.7 13.3 8.1 ;
        RECT 11.45 5.45 11.7 8.1 ;
        RECT 8.9 6.2 9.15 8.1 ;
        RECT 6.1 5.45 6.35 8.1 ;
        RECT 3.05 5.45 3.3 8.1 ;
        RECT 1.45 6.2 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 17.2 0.6 ;
        RECT 15.5 0 15.75 1.8 ;
        RECT 12.35 0 12.6 1.8 ;
        RECT 11.45 0 11.7 1.8 ;
        RECT 8.9 0 9.15 1.8 ;
        RECT 6.1 0 6.35 1.4 ;
        RECT 3.05 0 3.3 1.8 ;
        RECT 2.15 0 2.4 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 11.2 2.85 11.7 3.15 ;
      LAYER MET2 ;
        RECT 11.2 2.85 11.7 3.15 ;
        RECT 11.25 2.8 11.65 3.2 ;
      LAYER VIA12 ;
        RECT 11.32 2.87 11.58 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.55 3.5 4.05 3.8 ;
      LAYER MET2 ;
        RECT 3.55 3.45 4.05 3.85 ;
      LAYER VIA12 ;
        RECT 3.67 3.52 3.93 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.35 4.8 16.85 5.15 ;
        RECT 16.35 4.75 16.8 5.15 ;
        RECT 16.35 0.95 16.6 7.15 ;
      LAYER MET2 ;
        RECT 16.35 4.8 16.85 5.1 ;
        RECT 16.4 4.75 16.8 5.15 ;
      LAYER VIA12 ;
        RECT 16.47 4.82 16.73 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.65 4.15 16.1 4.45 ;
        RECT 15.75 2.05 16 4.45 ;
        RECT 14.65 2.05 16 2.3 ;
        RECT 14.65 4.15 14.9 7.15 ;
        RECT 14.65 0.95 14.9 2.3 ;
      LAYER MET2 ;
        RECT 15.6 4.15 16.1 4.45 ;
        RECT 15.65 4.1 16.05 4.5 ;
      LAYER VIA12 ;
        RECT 15.72 4.17 15.98 4.43 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.25 4.15 13.75 4.45 ;
        RECT 5.7 4.8 6.2 5.1 ;
        RECT 5.7 2.2 6.2 2.5 ;
        RECT 5.8 2.2 6.1 5.1 ;
        RECT 2.3 5.7 2.55 7.15 ;
        RECT 0.75 2.2 2.5 2.5 ;
        RECT 2.1 2.15 2.35 2.55 ;
        RECT 0.6 5.7 2.55 5.95 ;
        RECT 0.75 4.15 1.5 4.45 ;
        RECT 0.75 0.95 1 5.95 ;
        RECT 0.6 5.7 0.85 7.15 ;
      LAYER MET2 ;
        RECT 13.25 4.1 13.75 4.5 ;
        RECT 1.1 5.45 13.65 5.75 ;
        RECT 13.35 4.1 13.65 5.75 ;
        RECT 1 4.1 1.5 4.5 ;
        RECT 1.1 4.1 1.4 5.75 ;
        RECT 2 2.2 6.2 2.5 ;
        RECT 5.75 2.15 6.15 2.55 ;
        RECT 2 2.15 2.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.12 4.17 1.38 4.43 ;
        RECT 2.12 2.22 2.38 2.48 ;
        RECT 5.82 2.22 6.08 2.48 ;
        RECT 13.37 4.17 13.63 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 14.9 2.8 15.3 3.2 ;
      RECT 14.55 2.85 15.35 3.15 ;
      RECT 12.25 2.1 12.75 2.5 ;
      RECT 12.25 1.55 12.65 2.5 ;
      RECT 7.45 1.5 7.85 1.9 ;
      RECT 7.4 1.55 12.65 1.85 ;
      RECT 12.3 4.75 12.7 5.15 ;
      RECT 8.4 4.75 8.8 5.15 ;
      RECT 8.35 4.8 12.75 5.1 ;
      RECT 10.5 4.1 10.9 4.5 ;
      RECT 9.35 4.1 9.75 4.5 ;
      RECT 7.7 4.1 8.2 4.5 ;
      RECT 4.9 4.1 5.35 4.5 ;
      RECT 4.9 4.15 10.95 4.45 ;
      RECT 9.7 2.8 10.1 3.2 ;
      RECT 7.75 2.8 8.15 3.2 ;
      RECT 7.7 2.85 10.2 3.15 ;
      RECT 8.45 3.45 8.85 3.85 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 13.95 4.75 14.45 5.15 ;
      RECT 2 3.45 2.5 3.85 ;
    LAYER VIA12 ;
      RECT 14.97 2.87 15.23 3.13 ;
      RECT 14.07 4.82 14.33 5.08 ;
      RECT 12.37 2.17 12.63 2.43 ;
      RECT 12.37 4.82 12.63 5.08 ;
      RECT 10.57 4.17 10.83 4.43 ;
      RECT 9.77 2.87 10.03 3.13 ;
      RECT 9.42 4.17 9.68 4.43 ;
      RECT 8.52 3.52 8.78 3.78 ;
      RECT 8.47 4.82 8.73 5.08 ;
      RECT 7.82 2.87 8.08 3.13 ;
      RECT 7.82 4.17 8.08 4.43 ;
      RECT 7.52 1.57 7.78 1.83 ;
      RECT 5.02 4.17 5.28 4.43 ;
      RECT 2.12 3.52 2.38 3.78 ;
    LAYER MET1 ;
      RECT 14.05 2.85 14.35 5.2 ;
      RECT 12.35 4.7 12.65 5.2 ;
      RECT 12.35 4.8 14.35 5.1 ;
      RECT 13.75 2.85 15.35 3.15 ;
      RECT 13.75 0.95 14 3.15 ;
      RECT 13.9 6.2 14.15 7.15 ;
      RECT 12.2 6.2 12.45 7.15 ;
      RECT 12.2 6.2 14.15 6.45 ;
      RECT 10.6 0.95 10.85 7.15 ;
      RECT 10.55 1.7 10.85 5.6 ;
      RECT 10.55 4.15 10.9 4.45 ;
      RECT 9.75 4.75 10 7.15 ;
      RECT 9.75 4.75 10.3 5 ;
      RECT 10.05 3.55 10.3 5 ;
      RECT 9.75 2.75 10.05 3.8 ;
      RECT 9.75 0.95 10 3.8 ;
      RECT 8.35 4.8 8.85 5.1 ;
      RECT 8.45 3.5 8.75 5.1 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 7.15 4.15 8.2 4.45 ;
      RECT 7.15 2.15 7.45 4.45 ;
      RECT 7.05 2.15 7.55 2.45 ;
      RECT 7.5 5.95 7.75 7.15 ;
      RECT 6.6 5.95 7.75 6.2 ;
      RECT 6.6 3.45 6.85 6.2 ;
      RECT 6.55 1.6 6.8 3.7 ;
      RECT 6.55 1.6 7.9 1.85 ;
      RECT 7.5 1.55 7.9 1.85 ;
      RECT 7.5 0.95 7.75 1.85 ;
      RECT 4.25 4.15 5.4 4.45 ;
      RECT 5 2.2 5.3 4.45 ;
      RECT 4.9 2.2 5.4 2.5 ;
      RECT 4.7 4.95 4.95 7.15 ;
      RECT 3.05 4.95 4.95 5.2 ;
      RECT 3.05 2.25 3.3 5.2 ;
      RECT 2 3.5 3.3 3.8 ;
      RECT 3.05 2.25 4.05 2.5 ;
      RECT 3.65 1.55 4.05 2.5 ;
      RECT 3.65 1.55 4.95 1.8 ;
      RECT 4.7 0.95 4.95 1.8 ;
      RECT 12.25 2.15 12.75 2.45 ;
      RECT 9.3 4.15 9.8 4.45 ;
      RECT 7.7 2.85 8.2 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsr_1 0 0 ;
  SIZE 18.7 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 18.7 8.1 ;
        RECT 17.05 5.45 17.3 8.1 ;
        RECT 13.75 6.7 14 8.1 ;
        RECT 11.3 6.2 11.55 8.1 ;
        RECT 8.5 5.45 8.75 8.1 ;
        RECT 5.45 5.45 5.7 8.1 ;
        RECT 3.85 6.2 4.1 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 18.7 0.6 ;
        RECT 17.05 0 17.3 1.8 ;
        RECT 15.3 0 15.55 1.8 ;
        RECT 13.05 0 13.3 1.8 ;
        RECT 11.3 0 11.55 1.8 ;
        RECT 8.5 0 8.75 1.4 ;
        RECT 5.45 0 5.7 1.8 ;
        RECT 4.55 0 4.8 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 11.7 4.15 12.2 4.45 ;
        RECT 9.55 4.15 10.6 4.45 ;
        RECT 9.45 2.15 9.95 2.45 ;
        RECT 9.55 2.15 9.85 4.45 ;
        RECT 6.65 4.15 7.8 4.45 ;
        RECT 7.3 2.2 7.8 2.5 ;
        RECT 7.4 2.2 7.7 4.45 ;
      LAYER MET2 ;
        RECT 7.3 4.15 12.2 4.45 ;
        RECT 11.75 4.1 12.15 4.5 ;
        RECT 10.1 4.1 10.6 4.5 ;
        RECT 7.3 4.1 7.75 4.5 ;
      LAYER VIA12 ;
        RECT 7.42 4.17 7.68 4.43 ;
        RECT 10.22 4.17 10.48 4.43 ;
        RECT 11.82 4.17 12.08 4.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.95 3.5 6.45 3.8 ;
      LAYER MET2 ;
        RECT 5.95 3.45 6.45 3.85 ;
      LAYER VIA12 ;
        RECT 6.07 3.52 6.33 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 17.9 4.8 18.4 5.15 ;
        RECT 17.9 4.75 18.35 5.15 ;
        RECT 17.9 0.95 18.15 7.15 ;
      LAYER MET2 ;
        RECT 17.9 4.8 18.4 5.1 ;
        RECT 17.95 4.75 18.35 5.15 ;
      LAYER VIA12 ;
        RECT 18.02 4.82 18.28 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.2 4.15 17.65 4.45 ;
        RECT 17.3 2.05 17.55 4.45 ;
        RECT 16.2 2.05 17.55 2.3 ;
        RECT 16.2 4.15 16.45 7.15 ;
        RECT 16.2 0.95 16.45 2.3 ;
      LAYER MET2 ;
        RECT 17.15 4.15 17.65 4.45 ;
        RECT 17.2 4.1 17.6 4.5 ;
      LAYER VIA12 ;
        RECT 17.27 4.17 17.53 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.95 4.15 14.45 4.45 ;
        RECT 3.4 4.15 3.9 4.45 ;
      LAYER MET2 ;
        RECT 13.95 4.1 14.45 4.5 ;
        RECT 3.5 5.45 14.35 5.75 ;
        RECT 14.05 4.1 14.35 5.75 ;
        RECT 3.4 4.1 3.9 4.5 ;
        RECT 3.5 4.1 3.8 5.75 ;
      LAYER VIA12 ;
        RECT 3.52 4.17 3.78 4.43 ;
        RECT 14.07 4.17 14.33 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 16.45 2.8 16.85 3.2 ;
      RECT 16.1 2.85 16.9 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 14.85 2.1 15.45 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 14.85 0.9 15.15 2.5 ;
      RECT 2.75 0.9 15.15 1.2 ;
      RECT 12.95 2.1 13.45 2.5 ;
      RECT 12.95 1.55 13.35 2.5 ;
      RECT 9.85 1.5 10.25 1.9 ;
      RECT 9.8 1.55 13.35 1.85 ;
      RECT 13 4.75 13.4 5.15 ;
      RECT 10.8 4.75 11.2 5.15 ;
      RECT 10.75 4.8 13.45 5.1 ;
      RECT 12.1 2.8 12.5 3.2 ;
      RECT 10.15 2.8 10.55 3.2 ;
      RECT 10.1 2.85 12.6 3.15 ;
      RECT 10.85 3.45 11.25 3.85 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 8.15 2.15 8.55 2.55 ;
      RECT 4.4 2.15 4.9 2.55 ;
      RECT 4.4 2.2 8.6 2.5 ;
      RECT 15.35 4.75 15.85 5.15 ;
      RECT 4.4 3.45 4.9 3.85 ;
    LAYER VIA12 ;
      RECT 16.52 2.87 16.78 3.13 ;
      RECT 15.47 4.82 15.73 5.08 ;
      RECT 15.07 2.17 15.33 2.43 ;
      RECT 13.07 2.17 13.33 2.43 ;
      RECT 13.07 4.82 13.33 5.08 ;
      RECT 12.17 2.87 12.43 3.13 ;
      RECT 10.92 3.52 11.18 3.78 ;
      RECT 10.87 4.82 11.13 5.08 ;
      RECT 10.22 2.87 10.48 3.13 ;
      RECT 9.92 1.57 10.18 1.83 ;
      RECT 8.22 2.22 8.48 2.48 ;
      RECT 4.52 2.22 4.78 2.48 ;
      RECT 4.52 3.52 4.78 3.78 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 15.45 2.85 15.7 7.15 ;
      RECT 13.05 4.7 13.35 5.2 ;
      RECT 13.05 4.8 15.85 5.1 ;
      RECT 14.45 2.85 16.9 3.15 ;
      RECT 14.45 0.95 14.7 3.15 ;
      RECT 14.6 6.2 14.85 7.15 ;
      RECT 12.9 6.2 13.15 7.15 ;
      RECT 12.9 6.2 14.85 6.45 ;
      RECT 12.15 4.75 12.4 7.15 ;
      RECT 12.15 4.75 12.7 5 ;
      RECT 12.45 3.55 12.7 5 ;
      RECT 12.15 2.75 12.45 3.8 ;
      RECT 12.15 0.95 12.4 3.8 ;
      RECT 10.75 4.8 11.25 5.1 ;
      RECT 10.85 3.5 11.15 5.1 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 9.9 5.95 10.15 7.15 ;
      RECT 9 5.95 10.15 6.2 ;
      RECT 9 3.45 9.25 6.2 ;
      RECT 8.95 1.6 9.2 3.7 ;
      RECT 8.95 1.6 10.3 1.85 ;
      RECT 9.9 1.55 10.3 1.85 ;
      RECT 9.9 0.95 10.15 1.85 ;
      RECT 8.1 4.8 8.6 5.1 ;
      RECT 8.2 2.2 8.5 5.1 ;
      RECT 8.1 2.2 8.6 2.5 ;
      RECT 7.1 4.95 7.35 7.15 ;
      RECT 5.45 4.95 7.35 5.2 ;
      RECT 5.45 2.25 5.7 5.2 ;
      RECT 4.4 3.5 5.7 3.8 ;
      RECT 5.45 2.25 6.45 2.5 ;
      RECT 6.05 1.55 6.45 2.5 ;
      RECT 6.05 1.55 7.35 1.8 ;
      RECT 7.1 0.95 7.35 1.8 ;
      RECT 4.7 5.7 4.95 7.15 ;
      RECT 3 5.7 3.25 7.15 ;
      RECT 3 5.7 4.95 5.95 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 4.5 2.15 4.75 2.55 ;
      RECT 3.15 2.2 4.9 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 14.95 2.15 15.45 2.45 ;
      RECT 12.95 2.15 13.45 2.45 ;
      RECT 10.1 2.85 10.6 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsr_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsrn_1 0 0 ;
  SIZE 20.45 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 20.45 8.1 ;
        RECT 18.8 5.45 19.05 8.1 ;
        RECT 15.5 6.7 15.75 8.1 ;
        RECT 13.9 5.45 14.15 8.1 ;
        RECT 11.3 6.2 11.55 8.1 ;
        RECT 8.5 5.45 8.75 8.1 ;
        RECT 5.45 5.45 5.7 8.1 ;
        RECT 3.85 6.2 4.1 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 20.45 0.6 ;
        RECT 18.8 0 19.05 1.8 ;
        RECT 17.05 0 17.3 1.8 ;
        RECT 14.8 0 15.05 1.8 ;
        RECT 13.9 0 14.15 1.8 ;
        RECT 11.3 0 11.55 1.8 ;
        RECT 8.5 0 8.75 1.4 ;
        RECT 5.45 0 5.7 1.8 ;
        RECT 4.55 0 4.8 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 13.65 2.85 14.15 3.15 ;
      LAYER MET2 ;
        RECT 13.65 2.8 14.15 3.2 ;
      LAYER VIA12 ;
        RECT 13.77 2.87 14.03 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.95 3.5 6.45 3.8 ;
      LAYER MET2 ;
        RECT 5.95 3.45 6.45 3.85 ;
      LAYER VIA12 ;
        RECT 6.07 3.52 6.33 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 19.65 4.8 20.15 5.15 ;
        RECT 19.65 4.75 20.1 5.15 ;
        RECT 19.65 0.95 19.9 7.15 ;
      LAYER MET2 ;
        RECT 19.65 4.8 20.15 5.1 ;
        RECT 19.7 4.75 20.1 5.15 ;
      LAYER VIA12 ;
        RECT 19.77 4.82 20.03 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 17.95 4.15 19.4 4.45 ;
        RECT 19.05 2.05 19.3 4.45 ;
        RECT 17.95 2.05 19.3 2.3 ;
        RECT 17.95 4.15 18.2 7.15 ;
        RECT 17.95 0.95 18.2 2.3 ;
      LAYER MET2 ;
        RECT 18.9 4.15 19.4 4.45 ;
        RECT 18.95 4.1 19.35 4.5 ;
      LAYER VIA12 ;
        RECT 19.02 4.17 19.28 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.7 4.15 16.2 4.45 ;
        RECT 3.4 4.15 3.9 4.45 ;
      LAYER MET2 ;
        RECT 15.7 4.1 16.2 4.5 ;
        RECT 3.5 5.45 16.1 5.75 ;
        RECT 15.8 4.1 16.1 5.75 ;
        RECT 3.4 4.1 3.9 4.5 ;
        RECT 3.5 4.1 3.8 5.75 ;
      LAYER VIA12 ;
        RECT 3.52 4.17 3.78 4.43 ;
        RECT 15.82 4.17 16.08 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 18.2 2.8 18.6 3.2 ;
      RECT 17.85 2.85 18.65 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 16.6 2.1 17.2 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 16.6 0.9 16.9 2.5 ;
      RECT 2.75 0.9 16.9 1.2 ;
      RECT 14.7 2.1 15.2 2.5 ;
      RECT 14.7 1.55 15.1 2.5 ;
      RECT 9.85 1.5 10.25 1.9 ;
      RECT 9.8 1.55 15.1 1.85 ;
      RECT 14.75 4.75 15.15 5.15 ;
      RECT 10.8 4.75 11.2 5.15 ;
      RECT 10.75 4.8 15.2 5.1 ;
      RECT 12.95 4.1 13.4 4.5 ;
      RECT 11.75 4.1 12.15 4.5 ;
      RECT 10.1 4.1 10.6 4.5 ;
      RECT 7.3 4.1 7.75 4.5 ;
      RECT 7.3 4.15 13.4 4.45 ;
      RECT 12.1 2.8 12.5 3.2 ;
      RECT 10.15 2.8 10.55 3.2 ;
      RECT 10.1 2.85 12.6 3.15 ;
      RECT 10.85 3.45 11.25 3.85 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 8.15 2.15 8.55 2.55 ;
      RECT 4.4 2.15 4.9 2.55 ;
      RECT 4.4 2.2 8.6 2.5 ;
      RECT 17.1 4.75 17.6 5.15 ;
      RECT 4.4 3.45 4.9 3.85 ;
    LAYER VIA12 ;
      RECT 18.27 2.87 18.53 3.13 ;
      RECT 17.22 4.82 17.48 5.08 ;
      RECT 16.82 2.17 17.08 2.43 ;
      RECT 14.82 2.17 15.08 2.43 ;
      RECT 14.82 4.82 15.08 5.08 ;
      RECT 13.02 4.17 13.28 4.43 ;
      RECT 12.17 2.87 12.43 3.13 ;
      RECT 11.82 4.17 12.08 4.43 ;
      RECT 10.92 3.52 11.18 3.78 ;
      RECT 10.87 4.82 11.13 5.08 ;
      RECT 10.22 2.87 10.48 3.13 ;
      RECT 10.22 4.17 10.48 4.43 ;
      RECT 9.92 1.57 10.18 1.83 ;
      RECT 8.22 2.22 8.48 2.48 ;
      RECT 7.42 4.17 7.68 4.43 ;
      RECT 4.52 2.22 4.78 2.48 ;
      RECT 4.52 3.52 4.78 3.78 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 17.2 2.85 17.45 7.15 ;
      RECT 14.8 4.7 15.1 5.2 ;
      RECT 14.8 4.8 17.6 5.1 ;
      RECT 16.2 2.85 18.65 3.15 ;
      RECT 16.2 0.95 16.45 3.15 ;
      RECT 16.35 6.2 16.6 7.15 ;
      RECT 14.65 6.2 14.9 7.15 ;
      RECT 14.65 6.2 16.6 6.45 ;
      RECT 13.05 0.95 13.3 7.15 ;
      RECT 13 1.7 13.3 5.55 ;
      RECT 12.95 4.15 13.4 4.45 ;
      RECT 12.15 4.75 12.4 7.15 ;
      RECT 12.15 4.75 12.7 5 ;
      RECT 12.45 3.55 12.7 5 ;
      RECT 12.15 2.75 12.45 3.8 ;
      RECT 12.15 0.95 12.4 3.8 ;
      RECT 10.75 4.8 11.25 5.1 ;
      RECT 10.85 3.5 11.15 5.1 ;
      RECT 10.8 3.5 11.3 3.8 ;
      RECT 9.55 4.15 10.6 4.45 ;
      RECT 9.55 2.15 9.85 4.45 ;
      RECT 9.45 2.15 9.95 2.45 ;
      RECT 9.9 5.95 10.15 7.15 ;
      RECT 9 5.95 10.15 6.2 ;
      RECT 9 3.45 9.25 6.2 ;
      RECT 8.95 1.6 9.2 3.7 ;
      RECT 8.95 1.6 10.3 1.85 ;
      RECT 9.9 1.55 10.3 1.85 ;
      RECT 9.9 0.95 10.15 1.85 ;
      RECT 8.1 4.8 8.6 5.1 ;
      RECT 8.2 2.2 8.5 5.1 ;
      RECT 8.1 2.2 8.6 2.5 ;
      RECT 6.65 4.15 7.8 4.45 ;
      RECT 7.4 2.2 7.7 4.45 ;
      RECT 7.3 2.2 7.8 2.5 ;
      RECT 7.1 4.95 7.35 7.15 ;
      RECT 5.45 4.95 7.35 5.2 ;
      RECT 5.45 2.25 5.7 5.2 ;
      RECT 4.4 3.5 5.7 3.8 ;
      RECT 5.45 2.25 6.45 2.5 ;
      RECT 6.05 1.55 6.45 2.5 ;
      RECT 6.05 1.55 7.35 1.8 ;
      RECT 7.1 0.95 7.35 1.8 ;
      RECT 4.7 5.7 4.95 7.15 ;
      RECT 3 5.7 3.25 7.15 ;
      RECT 3 5.7 4.95 5.95 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 4.5 2.15 4.75 2.55 ;
      RECT 3.15 2.2 4.9 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 16.7 2.15 17.2 2.45 ;
      RECT 14.7 2.15 15.2 2.45 ;
      RECT 11.7 4.15 12.2 4.45 ;
      RECT 10.1 2.85 10.6 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsrn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dlat_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlat_1 0 0 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET2 ;
        RECT 5.2 4.1 5.7 4.5 ;
        RECT 3.45 4.15 5.7 4.45 ;
        RECT 3.5 4.1 3.9 4.5 ;
      LAYER MET1 ;
        RECT 5.2 4.15 5.7 4.45 ;
        RECT 3.45 4.15 3.95 4.45 ;
      LAYER VIA12 ;
        RECT 3.57 4.17 3.83 4.43 ;
        RECT 5.32 4.17 5.58 4.43 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 9 8.1 ;
        RECT 7.3 5.45 7.55 8.1 ;
        RECT 4.85 5.45 5.1 8.1 ;
        RECT 1.45 6.25 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9 0.6 ;
        RECT 7.3 0 7.55 1.8 ;
        RECT 4.7 0 5.1 1.8 ;
        RECT 1.45 0 1.85 1.8 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 1.85 4.1 2.35 4.5 ;
      LAYER MET1 ;
        RECT 1.85 4.15 2.35 4.45 ;
      LAYER VIA12 ;
        RECT 1.97 4.17 2.23 4.43 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET2 ;
        RECT 8.15 4.8 8.65 5.1 ;
        RECT 8.2 4.75 8.6 5.15 ;
      LAYER MET1 ;
        RECT 8.15 4.8 8.65 5.1 ;
        RECT 8.15 4.75 8.55 5.15 ;
        RECT 8.15 0.95 8.4 7.15 ;
      LAYER VIA12 ;
        RECT 8.27 4.82 8.53 5.08 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 6.75 3.45 7.25 3.85 ;
      RECT 4.55 3.45 4.95 3.85 ;
      RECT 0.35 3.45 0.85 3.85 ;
      RECT 0.35 3.5 7.25 3.8 ;
      RECT 6.5 4.75 6.9 5.15 ;
      RECT 6.45 4.8 6.95 5.1 ;
    LAYER VIA12 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.57 4.82 6.83 5.08 ;
      RECT 4.62 3.52 4.88 3.78 ;
      RECT 0.47 3.52 0.73 3.78 ;
    LAYER MET1 ;
      RECT 6.45 4.75 6.7 7.15 ;
      RECT 6.45 4.75 6.85 5.3 ;
      RECT 6.45 4.8 6.95 5.1 ;
      RECT 6.45 4.8 7.8 5.05 ;
      RECT 7.5 2.05 7.8 5.05 ;
      RECT 6.45 2.05 7.8 2.3 ;
      RECT 6.45 0.95 6.7 2.3 ;
      RECT 5.7 5.25 5.95 7.15 ;
      RECT 5.95 1.95 6.2 5.5 ;
      RECT 2.6 4.7 3.1 5 ;
      RECT 2.7 2.55 3 5 ;
      RECT 2.7 2.55 6.2 2.85 ;
      RECT 5.7 0.95 5.95 2.2 ;
      RECT 3.15 5.45 3.4 7.15 ;
      RECT 1.15 5.45 3.4 5.7 ;
      RECT 1.15 2.05 1.4 5.7 ;
      RECT 1.1 4.15 1.55 4.45 ;
      RECT 1.15 2.05 3.4 2.3 ;
      RECT 3.15 0.95 3.4 2.3 ;
      RECT 0.6 0.95 0.85 7.15 ;
      RECT 0.5 3.45 0.85 3.85 ;
      RECT 0.35 3.5 0.85 3.8 ;
      RECT 0.45 3.45 0.85 3.8 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.5 3.5 5 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlat_1

MACRO gf180mcu_osu_sc_gp12t3v3__dlatn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlatn_1 0 0 ;
  SIZE 10.7 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 10.7 8.1 ;
        RECT 9 5.45 9.25 8.1 ;
        RECT 7.4 5.45 7.65 8.1 ;
        RECT 4.85 5.45 5.1 8.1 ;
        RECT 1.45 6.25 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 10.7 0.6 ;
        RECT 9 0 9.25 1.8 ;
        RECT 7.4 0 7.65 1.8 ;
        RECT 4.7 0 5.1 1.8 ;
        RECT 1.45 0 1.85 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.05 2.55 7.55 2.85 ;
      LAYER MET2 ;
        RECT 7.05 2.5 7.55 2.9 ;
      LAYER VIA12 ;
        RECT 7.17 2.57 7.43 2.83 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 4.15 2.35 4.45 ;
      LAYER MET2 ;
        RECT 1.85 4.1 2.35 4.5 ;
      LAYER VIA12 ;
        RECT 1.97 4.17 2.23 4.43 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.85 4.8 10.35 5.1 ;
        RECT 9.85 4.75 10.25 5.15 ;
        RECT 9.85 0.95 10.1 7.15 ;
      LAYER MET2 ;
        RECT 9.85 4.8 10.35 5.1 ;
        RECT 9.9 4.75 10.3 5.15 ;
      LAYER VIA12 ;
        RECT 9.97 4.82 10.23 5.08 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 8.45 3.45 8.95 3.85 ;
      RECT 4.55 3.45 4.95 3.85 ;
      RECT 0.35 3.45 0.85 3.85 ;
      RECT 0.35 3.5 8.95 3.8 ;
      RECT 8.2 4.75 8.6 5.15 ;
      RECT 8.15 4.8 8.65 5.1 ;
      RECT 6.45 4.1 6.95 4.5 ;
      RECT 5.2 4.1 5.7 4.5 ;
      RECT 3.5 4.1 3.9 4.5 ;
      RECT 3.45 4.15 6.95 4.45 ;
    LAYER VIA12 ;
      RECT 8.57 3.52 8.83 3.78 ;
      RECT 8.27 4.82 8.53 5.08 ;
      RECT 6.57 4.17 6.83 4.43 ;
      RECT 5.32 4.17 5.58 4.43 ;
      RECT 4.62 3.52 4.88 3.78 ;
      RECT 3.57 4.17 3.83 4.43 ;
      RECT 0.47 3.52 0.73 3.78 ;
    LAYER MET1 ;
      RECT 8.15 4.75 8.4 7.15 ;
      RECT 8.15 4.75 8.55 5.3 ;
      RECT 8.15 4.8 8.65 5.1 ;
      RECT 8.15 4.8 9.5 5.05 ;
      RECT 9.2 2.05 9.5 5.05 ;
      RECT 8.15 2.05 9.5 2.3 ;
      RECT 8.15 0.95 8.4 2.3 ;
      RECT 6.55 0.95 6.8 7.15 ;
      RECT 6.55 4.1 6.95 4.5 ;
      RECT 6.45 4.15 6.95 4.45 ;
      RECT 5.7 5.25 5.95 7.15 ;
      RECT 5.95 1.95 6.2 5.5 ;
      RECT 2.6 4.7 3.1 5 ;
      RECT 2.7 2.55 3 5 ;
      RECT 2.7 2.55 6.2 2.85 ;
      RECT 5.7 0.95 5.95 2.2 ;
      RECT 3.15 5.45 3.4 7.15 ;
      RECT 1.15 5.45 3.4 5.7 ;
      RECT 1.15 2.05 1.4 5.7 ;
      RECT 1.1 4.15 1.55 4.45 ;
      RECT 1.15 2.05 3.4 2.3 ;
      RECT 3.15 0.95 3.4 2.3 ;
      RECT 0.6 0.95 0.85 7.15 ;
      RECT 0.5 3.45 0.85 3.85 ;
      RECT 0.35 3.5 0.85 3.8 ;
      RECT 0.45 3.45 0.85 3.8 ;
      RECT 8.45 3.5 8.95 3.8 ;
      RECT 5.2 4.15 5.7 4.45 ;
      RECT 4.5 3.5 5 3.8 ;
      RECT 3.45 4.15 3.95 4.45 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlatn_1

MACRO gf180mcu_osu_sc_gp12t3v3__fill_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_1 0 0 ;
  SIZE 0.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 0.1 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.1 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_1

MACRO gf180mcu_osu_sc_gp12t3v3__fill_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_16 0 0 ;
  SIZE 1.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 1.6 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 1.6 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_16

MACRO gf180mcu_osu_sc_gp12t3v3__fill_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_2 0 0 ;
  SIZE 0.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 0.2 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.2 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_2

MACRO gf180mcu_osu_sc_gp12t3v3__fill_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_4 0 0 ;
  SIZE 0.4 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 0.4 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.4 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_4

MACRO gf180mcu_osu_sc_gp12t3v3__fill_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_8 0 0 ;
  SIZE 0.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.8 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_8

MACRO gf180mcu_osu_sc_gp12t3v3__inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_1 0 0 ;
  SIZE 2.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.2 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_1

MACRO gf180mcu_osu_sc_gp12t3v3__inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_16 0 0 ;
  SIZE 15 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15 8.1 ;
        RECT 14.15 5.45 14.4 8.1 ;
        RECT 12.45 5.45 12.7 8.1 ;
        RECT 10.75 5.45 11 8.1 ;
        RECT 9.05 5.45 9.3 8.1 ;
        RECT 7.35 5.45 7.6 8.1 ;
        RECT 5.65 5.45 5.9 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15 0.6 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 12.45 0 12.7 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 9.05 0 9.3 1.8 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.3 0.95 13.55 7.15 ;
        RECT 1.4 4.45 13.55 4.7 ;
        RECT 13.15 4.1 13.55 4.7 ;
        RECT 1.4 2.05 13.55 2.3 ;
        RECT 11.6 0.95 11.85 7.15 ;
        RECT 9.9 0.95 10.15 7.15 ;
        RECT 8.2 0.95 8.45 7.15 ;
        RECT 6.5 0.95 6.75 7.15 ;
        RECT 4.8 0.95 5.05 7.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 13.15 4.1 13.65 4.5 ;
      LAYER VIA12 ;
        RECT 13.27 4.17 13.53 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_16

MACRO gf180mcu_osu_sc_gp12t3v3__inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_2 0 0 ;
  SIZE 3.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.2 8.1 ;
        RECT 2.3 5.45 2.55 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 3.5 1.15 3.8 ;
      LAYER MET2 ;
        RECT 0.65 3.45 1.15 3.85 ;
      LAYER VIA12 ;
        RECT 0.77 3.52 1.03 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 4.15 2 4.45 ;
        RECT 1.4 4 1.85 4.55 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 1.5 4.1 2 4.5 ;
      LAYER VIA12 ;
        RECT 1.62 4.17 1.88 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_2

MACRO gf180mcu_osu_sc_gp12t3v3__inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_4 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 4.45 3.35 4.7 ;
        RECT 2.95 4.1 3.35 4.7 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 2.95 4.1 3.45 4.5 ;
      LAYER VIA12 ;
        RECT 3.07 4.17 3.33 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_4

MACRO gf180mcu_osu_sc_gp12t3v3__inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_8 0 0 ;
  SIZE 8.15 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 8.15 8.1 ;
        RECT 7.35 5.45 7.6 8.1 ;
        RECT 5.65 5.45 5.9 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.15 0.6 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.5 0.95 6.75 7.15 ;
        RECT 1.4 4.45 6.75 4.7 ;
        RECT 6.35 4.1 6.75 4.7 ;
        RECT 1.4 2.05 6.75 2.3 ;
        RECT 4.8 0.95 5.05 7.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 6.35 4.1 6.85 4.5 ;
      LAYER VIA12 ;
        RECT 6.47 4.17 6.73 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_8

MACRO gf180mcu_osu_sc_gp12t3v3__lshifdown
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifdown 0 0 ;
  SIZE 5.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 2.9 7.5 5.2 8.1 ;
        RECT 3.45 5.45 3.75 8.1 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.3 8.1 ;
        RECT 0.55 5.45 0.85 8.1 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.2 0.6 ;
        RECT 3.45 0 3.75 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.3 4.15 4.7 4.45 ;
        RECT 4.35 0.95 4.65 7.15 ;
      LAYER MET2 ;
        RECT 4.25 4.1 4.75 4.5 ;
      LAYER VIA12 ;
        RECT 4.37 4.17 4.63 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 3.5 4.75 4 5.15 ;
      RECT 1.35 4.75 1.85 5.15 ;
      RECT 1.35 4.8 4 5.1 ;
    LAYER VIA12 ;
      RECT 3.62 4.82 3.88 5.08 ;
      RECT 1.47 4.82 1.73 5.08 ;
    LAYER MET1 ;
      RECT 1.45 0.95 1.75 7.15 ;
      RECT 1.35 4.8 1.85 5.1 ;
      RECT 3.5 4.8 4 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifdown

MACRO gf180mcu_osu_sc_gp12t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifup 0 0 ;
  SIZE 7.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.3 8.1 ;
        RECT 0.55 5.45 0.85 8.1 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.9 7.5 7.8 8.1 ;
        RECT 6.05 5.45 6.35 8.1 ;
        RECT 4.35 5.45 4.65 8.1 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 7.8 0.6 ;
        RECT 6.05 0 6.35 1.8 ;
        RECT 4.35 0 4.65 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4 2.2 4.5 2.5 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 4 2.15 4.5 2.55 ;
        RECT 0.6 2.2 4.5 2.5 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
        RECT 4.12 2.22 4.38 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.9 4.15 7.3 4.45 ;
        RECT 6.95 0.95 7.25 7.15 ;
      LAYER MET2 ;
        RECT 6.85 4.1 7.35 4.5 ;
      LAYER VIA12 ;
        RECT 6.97 4.17 7.23 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 6.1 4.75 6.6 5.15 ;
      RECT 4.55 4.75 4.95 5.15 ;
      RECT 4.5 4.8 6.6 5.1 ;
      RECT 4.5 2.85 5 3.25 ;
      RECT 1.35 2.85 1.85 3.25 ;
      RECT 1.35 2.9 5 3.2 ;
    LAYER VIA12 ;
      RECT 6.22 4.82 6.48 5.08 ;
      RECT 4.62 2.92 4.88 3.18 ;
      RECT 4.62 4.82 4.88 5.08 ;
      RECT 1.47 2.92 1.73 3.18 ;
    LAYER MET1 ;
      RECT 5.25 0.95 5.55 7.15 ;
      RECT 4.8 4 5.55 4.45 ;
      RECT 3.45 0.95 3.75 7.15 ;
      RECT 4.55 4.75 5 5.2 ;
      RECT 3.45 4.8 5 5.1 ;
      RECT 1.45 0.95 1.75 7.15 ;
      RECT 1.35 2.9 1.85 3.2 ;
      RECT 6.1 4.8 6.6 5.1 ;
      RECT 4.5 2.9 5 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifup

MACRO gf180mcu_osu_sc_gp12t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__mux2_1 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 3.45 2.85 3.85 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.75 4.1 4.25 4.5 ;
        RECT 3.95 0.95 4.2 7.15 ;
      LAYER MET2 ;
        RECT 3.75 4.1 4.25 4.5 ;
      LAYER VIA12 ;
        RECT 3.87 4.17 4.13 4.43 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.85 1.05 3.15 ;
      LAYER MET2 ;
        RECT 0.55 2.8 1.05 3.2 ;
      LAYER VIA12 ;
        RECT 0.67 2.87 0.93 3.13 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.75 3.5 5.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
      LAYER MET2 ;
        RECT 3 4.75 3.5 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 4.82 3.38 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.4 4.15 2 4.45 ;
      RECT 1.4 2.2 2 2.5 ;
  END
END gf180mcu_osu_sc_gp12t3v3__mux2_1

MACRO gf180mcu_osu_sc_gp12t3v3__nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nand2_1 0 0 ;
  SIZE 3.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.1 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.1 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 2.85 2.4 3.15 ;
      LAYER MET2 ;
        RECT 1.9 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.02 2.87 2.28 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 4.15 1.8 4.45 ;
        RECT 1.4 1.9 1.65 7.15 ;
        RECT 0.7 1.9 1.65 2.15 ;
        RECT 0.7 0.95 0.95 2.15 ;
      LAYER MET2 ;
        RECT 1.3 4.1 1.8 4.5 ;
      LAYER VIA12 ;
        RECT 1.42 4.17 1.68 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__nand2_1

MACRO gf180mcu_osu_sc_gp12t3v3__nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor2_1 0 0 ;
  SIZE 2.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.5 0.95 3.8 ;
      LAYER MET2 ;
        RECT 0.45 3.45 0.95 3.85 ;
      LAYER VIA12 ;
        RECT 0.57 3.52 0.83 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 4.75 2.2 7.15 ;
        RECT 1.25 4.75 2.2 5 ;
        RECT 1.15 4.15 1.65 4.45 ;
        RECT 1.25 0.95 1.5 5 ;
      LAYER MET2 ;
        RECT 1.15 4.1 1.65 4.5 ;
      LAYER VIA12 ;
        RECT 1.27 4.17 1.53 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__nor2_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai21_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 2.95 5.45 3.2 8.1 ;
        RECT 0.65 5.45 0.9 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 1.35 0 1.6 1.5 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.5 0.95 3.8 ;
      LAYER MET2 ;
        RECT 0.45 3.45 0.95 3.85 ;
      LAYER VIA12 ;
        RECT 0.57 3.52 0.83 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4.15 1.95 4.45 ;
      LAYER MET2 ;
        RECT 1.45 4.1 1.95 4.5 ;
      LAYER VIA12 ;
        RECT 1.57 4.17 1.83 4.43 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 3.5 2.7 3.8 ;
      LAYER MET2 ;
        RECT 2.2 3.45 2.7 3.85 ;
      LAYER VIA12 ;
        RECT 2.32 3.52 2.58 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 4.8 3.35 5.1 ;
        RECT 3.05 0.95 3.3 2.5 ;
        RECT 2.95 2.25 3.2 5.1 ;
        RECT 2.1 4.8 2.35 7.15 ;
      LAYER MET2 ;
        RECT 2.85 4.75 3.35 5.15 ;
      LAYER VIA12 ;
        RECT 2.97 4.82 3.23 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.75 2.45 2 ;
      RECT 2.2 0.95 2.45 2 ;
      RECT 0.5 0.95 0.75 2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai21_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai22_1 0 0 ;
  SIZE 5.3 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.3 8.1 ;
        RECT 3.5 5.45 3.75 8.1 ;
        RECT 0.65 5.45 0.9 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.3 0.6 ;
        RECT 1.35 0 1.6 1.6 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.5 0.95 3.8 ;
      LAYER MET2 ;
        RECT 0.45 3.45 0.95 3.85 ;
      LAYER VIA12 ;
        RECT 0.57 3.52 0.83 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4.15 1.95 4.45 ;
      LAYER MET2 ;
        RECT 1.45 4.1 1.95 4.5 ;
      LAYER VIA12 ;
        RECT 1.57 4.17 1.83 4.43 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 3.5 2.7 3.8 ;
      LAYER MET2 ;
        RECT 2.2 3.45 2.7 3.85 ;
      LAYER VIA12 ;
        RECT 2.32 3.52 2.58 3.78 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.15 3.5 3.65 3.8 ;
      LAYER MET2 ;
        RECT 3.15 3.45 3.65 3.85 ;
      LAYER VIA12 ;
        RECT 3.27 3.52 3.53 3.78 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.3 4.15 4.8 4.45 ;
        RECT 4.4 0.85 4.7 1.35 ;
        RECT 2.1 4.9 4.65 5.2 ;
        RECT 4.4 0.85 4.65 5.2 ;
        RECT 2.1 4.9 2.35 7.15 ;
        RECT 2.95 0.9 3.45 1.2 ;
        RECT 3.05 0.9 3.3 1.6 ;
      LAYER MET2 ;
        RECT 4.3 4.1 4.8 4.5 ;
        RECT 4.35 0.85 4.75 1.35 ;
        RECT 2.95 0.9 4.75 1.2 ;
        RECT 2.95 0.85 3.45 1.25 ;
      LAYER VIA12 ;
        RECT 3.07 0.92 3.33 1.18 ;
        RECT 4.42 4.17 4.68 4.43 ;
        RECT 4.42 0.97 4.68 1.23 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.85 4.15 2.1 ;
      RECT 3.9 0.95 4.15 2.1 ;
      RECT 2.2 0.95 2.45 2.1 ;
      RECT 0.5 0.95 0.75 2.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai22_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai31_1 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 3.85 5.45 4.1 8.1 ;
        RECT 1.05 5.45 1.3 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 2.25 0 2.5 1.5 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 2.85 1.45 3.15 ;
      LAYER MET2 ;
        RECT 0.95 2.8 1.45 3.2 ;
      LAYER VIA12 ;
        RECT 1.07 2.87 1.33 3.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 2.85 2.3 3.15 ;
      LAYER MET2 ;
        RECT 1.8 2.8 2.3 3.2 ;
      LAYER VIA12 ;
        RECT 1.92 2.87 2.18 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 4.15 3.05 4.45 ;
      LAYER MET2 ;
        RECT 2.55 4.1 3.05 4.5 ;
      LAYER VIA12 ;
        RECT 2.67 4.17 2.93 4.43 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 2.85 3.6 3.15 ;
      LAYER MET2 ;
        RECT 3.1 2.8 3.6 3.2 ;
      LAYER VIA12 ;
        RECT 3.22 2.87 3.48 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.8 4.25 5.1 ;
        RECT 3.95 0.95 4.2 2.5 ;
        RECT 3.85 2.25 4.1 5.1 ;
        RECT 3 4.8 3.25 7.15 ;
      LAYER MET2 ;
        RECT 3.75 4.75 4.25 5.15 ;
      LAYER VIA12 ;
        RECT 3.87 4.82 4.13 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.75 3.35 2 ;
      RECT 3.1 0.95 3.35 2 ;
      RECT 1.4 0.95 1.65 2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai31_1

MACRO gf180mcu_osu_sc_gp12t3v3__or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__or2_1 0 0 ;
  SIZE 3.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.8 8.1 ;
        RECT 1.95 5.45 2.35 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 3.5 1.4 3.8 ;
      LAYER MET2 ;
        RECT 0.9 3.45 1.4 3.85 ;
      LAYER VIA12 ;
        RECT 1.02 3.52 1.28 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.85 2.15 3.15 ;
      LAYER MET2 ;
        RECT 1.65 2.8 2.15 3.2 ;
      LAYER VIA12 ;
        RECT 1.77 2.87 2.03 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 4.8 3.45 5.1 ;
        RECT 2.95 0.95 3.2 7.15 ;
      LAYER MET2 ;
        RECT 2.95 4.75 3.45 5.15 ;
      LAYER VIA12 ;
        RECT 3.07 4.82 3.33 5.08 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.2 4.1 2.7 4.5 ;
    LAYER VIA12 ;
      RECT 2.32 4.17 2.58 4.43 ;
    LAYER MET1 ;
      RECT 0.55 5.25 0.8 7.15 ;
      RECT 0.4 2.2 0.65 5.5 ;
      RECT 0.4 4.15 2.7 4.45 ;
      RECT 0.4 2.2 1.5 2.45 ;
      RECT 1.25 0.95 1.5 2.45 ;
  END
END gf180mcu_osu_sc_gp12t3v3__or2_1

MACRO gf180mcu_osu_sc_gp12t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tbuf_1 0 0 ;
  SIZE 5.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.2 8.1 ;
        RECT 3.55 5.45 3.8 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.2 0.6 ;
        RECT 3.55 0 3.8 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 2.25 3.5 2.55 ;
      LAYER MET2 ;
        RECT 3 2.2 3.5 2.6 ;
      LAYER VIA12 ;
        RECT 3.12 2.27 3.38 2.53 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 5.45 3.05 7.15 ;
        RECT 1.95 1.55 3.05 1.8 ;
        RECT 2.8 0.95 3.05 1.8 ;
        RECT 2.45 3.5 2.95 3.8 ;
        RECT 1.95 4.25 2.8 4.5 ;
        RECT 2.55 2.75 2.8 4.5 ;
        RECT 1.95 5.45 3.05 5.7 ;
        RECT 1.95 2.75 2.8 3 ;
        RECT 1.95 4.25 2.2 5.7 ;
        RECT 1.95 1.55 2.2 3 ;
      LAYER MET2 ;
        RECT 2.45 3.45 2.95 3.85 ;
      LAYER VIA12 ;
        RECT 2.57 3.52 2.83 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 4.3 4.75 4.8 5.15 ;
      RECT 2.45 4.75 2.95 5.15 ;
      RECT 2.45 4.8 4.8 5.1 ;
    LAYER VIA12 ;
      RECT 4.42 4.82 4.68 5.08 ;
      RECT 2.57 4.82 2.83 5.08 ;
    LAYER MET1 ;
      RECT 4.4 0.95 4.65 7.15 ;
      RECT 4.3 4.8 4.8 5.1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 3.35 2 3.65 ;
      RECT 2.45 4.8 2.95 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tbuf_1

MACRO gf180mcu_osu_sc_gp12t3v3__tieh
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tieh 0 0 ;
  SIZE 2.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.2 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 4.8 1.8 5.1 ;
        RECT 1.4 4.75 1.65 7.15 ;
      LAYER MET2 ;
        RECT 1.3 4.75 1.8 5.15 ;
      LAYER VIA12 ;
        RECT 1.42 4.82 1.68 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.15 2.2 1.65 2.45 ;
      RECT 1.4 0.95 1.65 2.45 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tieh

MACRO gf180mcu_osu_sc_gp12t3v3__tiel
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tiel 0 0 ;
  SIZE 2.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.2 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 2.1 1.8 2.4 ;
        RECT 1.4 0.95 1.65 2.45 ;
      LAYER MET2 ;
        RECT 1.3 2.05 1.8 2.45 ;
      LAYER VIA12 ;
        RECT 1.42 2.12 1.68 2.38 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 4.85 1.65 7.15 ;
      RECT 1.15 4.85 1.65 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tiel

MACRO gf180mcu_osu_sc_gp12t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tinv_1 0 0 ;
  SIZE 3.65 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.65 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.65 0.6 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4.8 1.95 5.1 ;
      LAYER MET2 ;
        RECT 1.45 4.75 1.95 5.15 ;
      LAYER VIA12 ;
        RECT 1.57 4.82 1.83 5.08 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.7 2.2 3.2 2.5 ;
        RECT 1 2.2 1.5 2.5 ;
      LAYER MET2 ;
        RECT 2.7 2.15 3.2 2.55 ;
        RECT 1 2.2 3.2 2.5 ;
        RECT 1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.12 2.22 1.38 2.48 ;
        RECT 2.82 2.22 3.08 2.48 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 5.45 3.05 7.15 ;
        RECT 2.2 1.55 3.05 1.8 ;
        RECT 2.8 0.95 3.05 1.8 ;
        RECT 2.2 5.45 3.05 5.7 ;
        RECT 2.05 3.5 2.6 3.8 ;
        RECT 2.2 1.55 2.45 5.7 ;
      LAYER MET2 ;
        RECT 2.05 3.45 2.55 3.85 ;
      LAYER VIA12 ;
        RECT 2.17 3.52 2.43 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.7 4.75 3.2 5.15 ;
      RECT 2.8 4.15 3.1 5.15 ;
      RECT 0.35 4.1 0.85 4.5 ;
      RECT 0.35 4.15 3.1 4.45 ;
    LAYER VIA12 ;
      RECT 2.82 4.82 3.08 5.08 ;
      RECT 0.47 4.17 0.73 4.43 ;
    LAYER MET1 ;
      RECT 0.55 5.45 0.8 7.15 ;
      RECT 0.5 1.8 0.75 5.7 ;
      RECT 0.35 4.15 0.85 4.45 ;
      RECT 0.55 0.95 0.8 2.05 ;
      RECT 2.7 4.8 3.2 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tinv_1

MACRO gf180mcu_osu_sc_gp12t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xnor2_1 0 0 ;
  SIZE 6.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 6.2 8.1 ;
        RECT 4.5 5.45 4.75 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.2 0.6 ;
        RECT 4.5 0 4.75 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.55 3.5 4.05 3.8 ;
        RECT 1.25 2.2 1.75 2.5 ;
      LAYER MET2 ;
        RECT 3.6 3.45 4 3.85 ;
        RECT 3.65 0.9 3.95 3.9 ;
        RECT 1.35 0.9 3.95 1.2 ;
        RECT 1.3 2.15 1.7 2.55 ;
        RECT 1.35 0.9 1.65 2.6 ;
      LAYER VIA12 ;
        RECT 1.37 2.22 1.63 2.48 ;
        RECT 3.67 3.52 3.93 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.35 2.2 4.85 2.5 ;
      LAYER MET2 ;
        RECT 4.35 2.2 4.85 2.5 ;
        RECT 4.4 2.15 4.8 2.55 ;
        RECT 4.45 2.1 4.75 2.6 ;
      LAYER VIA12 ;
        RECT 4.47 2.22 4.73 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 1.4 3.2 1.95 ;
        RECT 2.95 0.95 3.2 1.95 ;
        RECT 2.95 5.3 3.2 7.15 ;
        RECT 2.9 5.3 3.2 5.85 ;
      LAYER MET2 ;
        RECT 2.8 1.5 3.3 1.9 ;
        RECT 2.85 5.4 3.25 5.8 ;
        RECT 2.9 1.5 3.2 5.95 ;
      LAYER VIA12 ;
        RECT 2.92 5.47 3.18 5.73 ;
        RECT 2.92 1.57 3.18 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.35 0.95 5.6 7.15 ;
      RECT 2.55 4.15 5.6 4.45 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 3.5 3.3 3.8 ;
      RECT 3 2.2 3.3 3.8 ;
      RECT 2.9 2.2 3.4 2.5 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xnor2_1

MACRO gf180mcu_osu_sc_gp12t3v3__xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xor2_1 0 0 ;
  SIZE 6.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 6.2 8.1 ;
        RECT 4.5 5.45 4.75 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.2 0.6 ;
        RECT 4.5 0 4.75 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.25 2.2 1.75 2.5 ;
      LAYER MET2 ;
        RECT 1.25 2.2 1.75 2.5 ;
        RECT 1.3 2.15 1.7 2.55 ;
      LAYER VIA12 ;
        RECT 1.37 2.22 1.63 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 3.5 5.1 3.8 ;
      LAYER MET2 ;
        RECT 4.6 3.5 5.1 3.8 ;
        RECT 4.65 3.45 5.05 3.85 ;
        RECT 1.95 3.5 2.45 3.8 ;
        RECT 2 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.07 3.52 2.33 3.78 ;
        RECT 4.72 3.52 4.98 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 1.4 3.2 1.95 ;
        RECT 2.95 0.95 3.2 1.95 ;
        RECT 2.95 5.35 3.2 7.15 ;
        RECT 2.9 5.35 3.2 5.85 ;
      LAYER MET2 ;
        RECT 2.8 1.5 3.3 1.9 ;
        RECT 2.85 5.4 3.25 5.8 ;
        RECT 2.9 1.5 3.2 5.95 ;
      LAYER VIA12 ;
        RECT 2.92 5.47 3.18 5.73 ;
        RECT 2.92 1.57 3.18 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.35 0.95 5.6 7.15 ;
      RECT 2.55 4.8 5.6 5.1 ;
      RECT 4.05 2.2 5.6 2.5 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 4.15 4.05 4.45 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xor2_1

END LIBRARY
