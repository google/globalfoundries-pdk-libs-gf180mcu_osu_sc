* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffr_1 D Q QN CLK RN VDD VSS
X0 VDD a_41_109# a_145_109# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_173_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 a_122_14# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_122_14# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 VDD a_205_68# a_201_109# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_62_98# CLK a_112_109# VDD pmos_3p3 w=1.7u l=0.3u
X6 a_145_109# a_122_14# a_62_98# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_145_19# CLK a_62_98# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 a_62_98# a_122_14# a_112_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_112_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_205_68# a_184_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 VDD a_205_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X15 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X16 a_201_19# a_122_14# a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X17 VSS a_205_68# a_201_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X19 a_205_68# a_25_19# a_273_109# VDD pmos_3p3 w=1.7u l=0.3u
X20 a_273_109# a_184_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X21 VSS a_205_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X22 VSS a_62_98# a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD a_62_98# a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_112_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 VSS a_25_19# a_205_68# VSS nmos_3p3 w=0.85u l=0.3u
X26 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_173_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X28 a_201_109# CLK a_184_19# VDD pmos_3p3 w=1.7u l=0.3u
X29 a_184_19# a_122_14# a_173_109# VDD pmos_3p3 w=1.7u l=0.3u
X30 VSS a_41_109# a_145_19# VSS nmos_3p3 w=0.85u l=0.3u
X31 a_184_19# CLK a_173_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
