# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xnor2_1 0 0 ;
  SIZE 6.4 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 6.4 6.35 ;
        RECT 4.7 4.7 4.95 6.35 ;
        RECT 1.4 4.7 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 6.4 0.7 ;
        RECT 4.7 0 4.95 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.5 3.1 4 3.4 ;
        RECT 1.25 2.3 1.75 2.6 ;
      LAYER Metal2 ;
        RECT 3.55 3.05 4 3.45 ;
        RECT 3.7 1 4 3.45 ;
        RECT 3.6 3 3.95 3.5 ;
        RECT 1.35 1 4 1.3 ;
        RECT 1.3 2.25 1.7 2.65 ;
        RECT 1.35 1 1.65 2.7 ;
      LAYER Via1 ;
        RECT 1.37 2.32 1.63 2.58 ;
        RECT 3.62 3.12 3.88 3.38 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.55 2.3 5.05 2.6 ;
      LAYER Metal2 ;
        RECT 4.55 2.3 5.05 2.6 ;
        RECT 4.6 2.25 5 2.65 ;
        RECT 4.65 2.2 4.95 2.7 ;
      LAYER Via1 ;
        RECT 4.67 2.32 4.93 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 1.5 3.3 2.05 ;
        RECT 3.05 1.05 3.3 2.05 ;
        RECT 3.05 4.15 3.3 5.3 ;
        RECT 3 4.15 3.3 4.85 ;
      LAYER Metal2 ;
        RECT 2.9 1.6 3.4 2 ;
        RECT 2.95 4.2 3.35 4.6 ;
        RECT 3 4.15 3.3 4.85 ;
        RECT 2.95 1.6 3.25 4.6 ;
      LAYER Via1 ;
        RECT 3.02 4.27 3.28 4.53 ;
        RECT 3.02 1.67 3.28 1.93 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5.55 1.05 5.8 5.3 ;
      RECT 2.75 3.65 5.8 3.9 ;
      RECT 2.75 3 3.05 3.9 ;
      RECT 0.55 1.05 0.8 5.3 ;
      RECT 0.55 3.1 2.4 3.4 ;
      RECT 2.1 2.3 2.4 3.4 ;
      RECT 2.1 2.3 3.5 2.6 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xnor2_1
