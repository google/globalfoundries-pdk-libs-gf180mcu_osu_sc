* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dlat_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dlat_1 D Q CLK VDD VSS
X0 VDD a_10_19# a_77_70# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_52_58# CLK VSS VSS nmos_3p3 w=0.85u l=0.3u
X2 VDD a_20_14# a_10_19# VDD pmos_3p3 w=1.7u l=0.3u
X3 Q a_137_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_52_58# CLK VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 a_46_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_20_14# CLK a_46_19# VSS nmos_3p3 w=0.85u l=0.3u
X7 a_20_14# a_52_58# a_43_70# VDD pmos_3p3 w=1.7u l=0.3u
X8 VSS a_10_19# a_137_19# VSS nmos_3p3 w=0.85u l=0.3u
X9 VDD a_10_19# a_137_19# VDD pmos_3p3 w=1.7u l=0.3u
X10 a_77_19# a_52_58# a_20_14# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_77_70# CLK a_20_14# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_20_14# a_10_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 Q a_137_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 a_43_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS a_10_19# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
