# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xnor2_1 0 0 ;
  SIZE 6.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 6.2 8.3 ;
        RECT 4.5 5.55 4.75 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 6.2 0.7 ;
        RECT 4.5 0 4.75 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 3.6 4.05 3.9 ;
        RECT 1.25 2.3 1.75 2.6 ;
      LAYER Metal2 ;
        RECT 3.6 3.55 4 3.95 ;
        RECT 3.65 1 3.95 4 ;
        RECT 1.35 1 3.95 1.3 ;
        RECT 1.3 2.25 1.7 2.65 ;
        RECT 1.35 1 1.65 2.7 ;
      LAYER Via1 ;
        RECT 1.37 2.32 1.63 2.58 ;
        RECT 3.67 3.62 3.93 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.35 2.3 4.85 2.6 ;
      LAYER Metal2 ;
        RECT 4.35 2.3 4.85 2.6 ;
        RECT 4.4 2.25 4.8 2.65 ;
        RECT 4.45 2.2 4.75 2.7 ;
      LAYER Via1 ;
        RECT 4.47 2.32 4.73 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 1.5 3.2 2.05 ;
        RECT 2.95 1.05 3.2 2.05 ;
        RECT 2.95 5.4 3.2 7.25 ;
        RECT 2.9 5.4 3.2 5.95 ;
      LAYER Metal2 ;
        RECT 2.8 1.6 3.3 2 ;
        RECT 2.85 5.5 3.25 5.9 ;
        RECT 2.9 1.6 3.2 6.05 ;
      LAYER Via1 ;
        RECT 2.92 5.57 3.18 5.83 ;
        RECT 2.92 1.67 3.18 1.93 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5.35 1.05 5.6 7.25 ;
      RECT 2.55 4.25 5.6 4.55 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3.6 3.3 3.9 ;
      RECT 3 2.3 3.3 3.9 ;
      RECT 2.9 2.3 3.4 2.6 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xnor2_1
