magic
tech gf180mcuC
timestamp 1661874533
<< nwell >>
rect 0 61 78 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 53 19 59 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 53 70 59 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 34 53 36
rect 42 21 45 34
rect 50 21 53 34
rect 42 19 53 21
rect 59 34 69 36
rect 59 21 62 34
rect 67 21 69 34
rect 59 19 69 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 36 104
rect 25 72 28 102
rect 33 72 36 102
rect 25 70 36 72
rect 42 102 53 104
rect 42 77 45 102
rect 50 77 53 102
rect 42 70 53 77
rect 59 102 69 104
rect 59 72 62 102
rect 67 72 69 102
rect 59 70 69 72
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 45 21 50 34
rect 62 21 67 34
<< pdiffc >>
rect 11 72 16 102
rect 28 72 33 102
rect 45 77 50 102
rect 62 72 67 102
<< psubdiff >>
rect 9 10 19 12
rect 9 5 11 10
rect 16 5 19 10
rect 9 3 19 5
rect 33 10 43 12
rect 33 5 35 10
rect 40 5 43 10
rect 33 3 43 5
rect 57 10 67 12
rect 57 5 59 10
rect 64 5 67 10
rect 57 3 67 5
<< nsubdiff >>
rect 9 118 19 120
rect 9 113 11 118
rect 16 113 19 118
rect 9 111 19 113
rect 33 118 43 120
rect 33 113 35 118
rect 40 113 43 118
rect 33 111 43 113
rect 57 118 67 120
rect 57 113 59 118
rect 64 113 67 118
rect 57 111 67 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 53 104 59 109
rect 19 52 25 70
rect 36 68 42 70
rect 53 68 59 70
rect 36 67 59 68
rect 30 65 59 67
rect 30 59 32 65
rect 38 62 59 65
rect 38 59 42 62
rect 30 57 42 59
rect 19 50 31 52
rect 19 44 23 50
rect 29 44 31 50
rect 19 42 31 44
rect 36 44 42 57
rect 19 36 25 42
rect 36 38 59 44
rect 36 36 42 38
rect 53 36 59 38
rect 19 14 25 19
rect 36 14 42 19
rect 53 14 59 19
<< polycontact >>
rect 32 59 38 65
rect 23 44 29 50
<< metal1 >>
rect 0 118 78 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 78 118
rect 0 111 78 112
rect 11 102 16 104
rect 11 65 16 72
rect 28 102 33 111
rect 45 102 50 104
rect 45 76 50 77
rect 62 102 67 111
rect 28 70 33 72
rect 43 70 45 76
rect 51 70 53 76
rect 62 70 67 72
rect 11 59 32 65
rect 38 59 40 65
rect 11 34 16 59
rect 21 44 23 50
rect 29 44 31 50
rect 11 19 16 21
rect 28 34 33 36
rect 28 12 33 21
rect 45 34 50 70
rect 45 19 50 21
rect 62 34 67 36
rect 62 12 67 21
rect 0 11 78 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 78 11
rect 0 0 78 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 45 70 51 76
rect 23 44 29 50
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 43 76 53 77
rect 43 70 45 76
rect 51 70 53 76
rect 43 69 53 70
rect 22 50 30 51
rect 21 44 23 50
rect 29 44 31 50
rect 22 43 30 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 26 47 26 47 1 A
port 1 n
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 48 73 48 73 1 Y
port 2 n
<< end >>
