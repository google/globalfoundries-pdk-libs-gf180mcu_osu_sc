* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_and2_1 A B Y
X0 Y a_12_16 VDD VDD pmos_3p3 w=34 l=6
X1 VDD B a_12_16 VDD pmos_3p3 w=34 l=6
X2 a_12_16 A VDD VDD pmos_3p3 w=34 l=6
X3 Y a_12_16 GND GND nmos_3p3 w=17 l=6
X4 a_28_16 A a_12_16 GND nmos_3p3 w=17 l=6
X5 GND B a_28_16 GND nmos_3p3 w=17 l=6
.ends

