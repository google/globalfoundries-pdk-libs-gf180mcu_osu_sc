* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dff_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dff_1 D Q QN CLK VDD VSS
X0 a_19_16# CLK a_42_72# VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_161_44# QN VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS a_9_21# a_86_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_19_16# a_53_40# a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS a_161_44# QN VSS nfet_03p3 w=0.85u l=0.3u
X5 VDD a_19_16# a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X6 a_53_40# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 VSS a_19_16# a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_53_40# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 a_148_72# CLK a_125_21# VDD pfet_03p3 w=1.7u l=0.3u
X10 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X11 a_114_72# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X12 a_161_44# a_125_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 a_148_21# a_53_40# a_125_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X15 a_42_72# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 a_125_21# a_53_40# a_114_72# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_114_21# a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X18 a_161_44# a_125_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X19 a_86_72# a_53_40# a_19_16# VDD pfet_03p3 w=1.7u l=0.3u
X20 VDD a_161_44# a_148_72# VDD pfet_03p3 w=1.7u l=0.3u
X21 a_42_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 a_125_21# CLK a_114_21# VSS nfet_03p3 w=0.85u l=0.3u
X23 VDD a_9_21# a_86_72# VDD pfet_03p3 w=1.7u l=0.3u
X24 a_86_21# CLK a_19_16# VSS nfet_03p3 w=0.85u l=0.3u
X25 VSS a_161_44# a_148_21# VSS nfet_03p3 w=0.85u l=0.3u
.ends
