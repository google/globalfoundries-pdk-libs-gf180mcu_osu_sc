* NGSPICE file created from gf180mcu_osu_sc_9T_xnor2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_42_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_49_14# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_49_14# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 GND A a_9_19# GND nmos_3p3 w=0.85u l=0.3u
X4 VDD A a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_78_19# a_9_19# Y GND nmos_3p3 w=0.85u l=0.3u
X6 GND B a_78_19# GND nmos_3p3 w=0.85u l=0.3u
X7 a_78_70# A Y VDD pmos_3p3 w=1.7u l=0.3u
X8 a_42_19# A GND GND nmos_3p3 w=0.85u l=0.3u
X9 VDD B a_78_70# VDD pmos_3p3 w=1.7u l=0.3u
X10 Y a_49_14# a_42_19# GND nmos_3p3 w=0.85u l=0.3u
X11 a_49_14# B GND GND nmos_3p3 w=0.85u l=0.3u
