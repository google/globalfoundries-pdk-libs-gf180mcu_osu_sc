magic
tech gf180mcuC
timestamp 1661875326
<< nwell >>
rect 0 61 102 123
<< nmos >>
rect 19 19 25 36
rect 53 19 59 36
rect 73 19 79 36
<< pmos >>
rect 19 70 25 104
rect 53 70 59 104
rect 73 70 79 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 35 36
rect 25 21 28 34
rect 33 21 35 34
rect 25 19 35 21
rect 43 34 53 36
rect 43 21 45 34
rect 50 21 53 34
rect 43 19 53 21
rect 59 34 73 36
rect 59 21 62 34
rect 67 21 73 34
rect 59 19 73 21
rect 79 34 92 36
rect 79 21 85 34
rect 90 21 92 34
rect 79 19 92 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 35 104
rect 25 72 28 102
rect 33 72 35 102
rect 25 70 35 72
rect 43 102 53 104
rect 43 72 45 102
rect 50 72 53 102
rect 43 70 53 72
rect 59 102 73 104
rect 59 95 62 102
rect 67 95 73 102
rect 59 70 73 95
rect 79 102 92 104
rect 79 72 85 102
rect 90 72 92 102
rect 79 70 92 72
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 45 21 50 34
rect 62 21 67 34
rect 85 21 90 34
<< pdiffc >>
rect 11 72 16 102
rect 28 72 33 102
rect 45 72 50 102
rect 62 95 67 102
rect 85 72 90 102
<< psubdiff >>
rect 9 10 19 12
rect 9 5 11 10
rect 16 5 19 10
rect 9 3 19 5
rect 33 10 43 12
rect 33 5 35 10
rect 40 5 43 10
rect 33 3 43 5
rect 57 10 67 12
rect 57 5 59 10
rect 64 5 67 10
rect 57 3 67 5
rect 81 10 91 12
rect 81 5 83 10
rect 88 5 91 10
rect 81 3 91 5
<< nsubdiff >>
rect 9 118 19 120
rect 9 113 11 118
rect 16 113 19 118
rect 9 111 19 113
rect 33 118 43 120
rect 33 113 35 118
rect 40 113 43 118
rect 33 111 43 113
rect 57 118 67 120
rect 57 113 59 118
rect 64 113 67 118
rect 57 111 67 113
rect 81 118 91 120
rect 81 113 83 118
rect 88 113 91 118
rect 81 111 91 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
<< polysilicon >>
rect 19 104 25 109
rect 53 104 59 109
rect 73 104 79 109
rect 19 65 25 70
rect 12 62 25 65
rect 12 57 14 62
rect 19 58 25 62
rect 53 58 59 70
rect 73 68 79 70
rect 71 66 81 68
rect 71 61 73 66
rect 79 61 81 66
rect 71 59 81 61
rect 19 57 66 58
rect 12 55 66 57
rect 19 54 66 55
rect 19 53 79 54
rect 19 36 25 53
rect 61 49 79 53
rect 30 46 40 48
rect 30 40 32 46
rect 38 44 40 46
rect 38 40 59 44
rect 30 39 59 40
rect 30 38 40 39
rect 53 36 59 39
rect 73 36 79 49
rect 19 14 25 19
rect 53 14 59 19
rect 73 14 79 19
<< polycontact >>
rect 14 57 19 62
rect 73 61 79 66
rect 32 40 38 46
<< metal1 >>
rect 0 118 102 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 102 118
rect 0 111 102 112
rect 11 102 16 111
rect 11 70 16 72
rect 28 102 33 104
rect 28 67 33 72
rect 45 102 50 104
rect 11 57 13 63
rect 19 57 21 63
rect 28 61 31 67
rect 37 61 39 67
rect 28 46 33 61
rect 45 51 50 72
rect 62 102 67 104
rect 62 91 67 95
rect 85 102 90 104
rect 62 89 68 91
rect 62 81 68 83
rect 45 50 57 51
rect 28 40 32 46
rect 38 40 40 46
rect 45 44 49 50
rect 55 44 57 50
rect 45 43 57 44
rect 11 34 16 36
rect 11 12 16 21
rect 28 34 33 40
rect 28 19 33 21
rect 45 34 50 43
rect 45 19 50 21
rect 62 34 67 81
rect 73 67 79 69
rect 73 58 79 61
rect 62 19 67 21
rect 85 51 90 72
rect 85 50 95 51
rect 85 44 87 50
rect 93 44 95 50
rect 85 43 95 44
rect 85 34 90 43
rect 85 19 90 21
rect 0 11 102 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 102 11
rect 0 0 102 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 13 62 19 63
rect 13 57 14 62
rect 14 57 19 62
rect 31 61 37 67
rect 62 83 68 89
rect 49 44 55 50
rect 73 66 79 67
rect 73 61 79 66
rect 87 44 93 50
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 60 89 70 90
rect 60 83 62 89
rect 68 83 70 89
rect 60 82 70 83
rect 29 67 39 68
rect 71 67 81 68
rect 11 63 21 64
rect 11 57 13 63
rect 19 57 21 63
rect 29 61 31 67
rect 37 61 73 67
rect 79 61 81 67
rect 29 60 39 61
rect 71 60 81 61
rect 11 56 21 57
rect 47 50 57 51
rect 47 44 49 50
rect 55 44 57 50
rect 47 43 57 44
rect 85 50 95 51
rect 85 44 87 50
rect 93 44 95 50
rect 85 43 95 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 52 47 52 47 1 A
port 4 n
rlabel metal2 90 47 90 47 1 B
port 5 n
rlabel metal2 16 60 16 60 1 Sel
port 3 n
rlabel metal2 65 86 65 86 1 Y
port 2 n
<< end >>
