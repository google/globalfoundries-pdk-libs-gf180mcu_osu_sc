* NGSPICE file created from gf180mcu_osu_sc_12T_oai21_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y B a_8_16# GND nmos_3p3 w=0.85u l=0.3u
X1 GND A0 a_8_16# GND nmos_3p3 w=0.85u l=0.3u
X2 a_27_106# A0 VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD B Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y A1 a_27_106# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_8_16# A1 GND GND nmos_3p3 w=0.85u l=0.3u
