# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_tinv_1 0 0 ;
  SIZE 3.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.5 6.15 ;
        RECT 1.15 3.5 1.4 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.5 0.6 ;
        RECT 1.15 0 1.4 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 2.1 2.45 2.6 ;
      LAYER MET2 ;
        RECT 2.05 2.15 2.55 2.55 ;
      LAYER VIA12 ;
        RECT 2.17 2.22 2.43 2.48 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.5 2.2 1 2.5 ;
      LAYER MET2 ;
        RECT 0.5 2.15 1 2.55 ;
      LAYER VIA12 ;
        RECT 0.62 2.22 0.88 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.2 2.85 1.7 3.15 ;
      LAYER MET2 ;
        RECT 1.2 2.8 1.7 3.2 ;
      LAYER VIA12 ;
        RECT 1.32 2.87 1.58 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.45 3.5 2.95 3.8 ;
        RECT 2.7 1.55 2.95 3.8 ;
        RECT 2.55 3.4 2.8 5.2 ;
        RECT 2.55 0.95 2.8 1.8 ;
      LAYER MET2 ;
        RECT 2.45 3.45 2.95 3.85 ;
      LAYER VIA12 ;
        RECT 2.57 3.52 2.83 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_9T_tinv_1
