* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__nfet_01v8_lvt.0 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.44292+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.45748
+ k2 = {-0.040708+sky130_fd_pr__nfet_01v8_lvt__k2_diff_0}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {84096+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_0}
+ ua = {-1.5106e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_0}
+ ub = {2.3749e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_0}
+ uc = 4.4533e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_0}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.026527+sky130_fd_pr__nfet_01v8_lvt__u0_diff_0}
+ a0 = {1.5497+sky130_fd_pr__nfet_01v8_lvt__a0_diff_0}
+ keta = {-0.11251+sky130_fd_pr__nfet_01v8_lvt__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.8405+sky130_fd_pr__nfet_01v8_lvt__ags_diff_0}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_0}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11515019+sky130_fd_pr__nfet_01v8_lvt__voff_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.0396987+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_0}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.00043348+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_0}
+ etab = -0.00047191
+ dsub = 0.57273167
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.21192+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_0}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.014693
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.7058626e-5
+ alpha1 = 0.0
+ beta0 = 20.772941
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26953+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_0}
+ kt2 = -0.022714
+ at = 78553.0
+ ute = -1.0929
+ ua1 = 1.9956e-9
+ ub1 = -1.7256e-18
+ uc1 = -4.9957e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.1 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43904+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.45793
+ k2 = {-0.03517+sky130_fd_pr__nfet_01v8_lvt__k2_diff_1}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {42698+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_1}
+ ua = {-1.1127e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_1}
+ ub = {2.2971e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_1}
+ uc = 5.1465e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_1}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.032411+sky130_fd_pr__nfet_01v8_lvt__u0_diff_1}
+ a0 = {1.9169+sky130_fd_pr__nfet_01v8_lvt__a0_diff_1}
+ keta = {-0.18123+sky130_fd_pr__nfet_01v8_lvt__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.5934+sky130_fd_pr__nfet_01v8_lvt__ags_diff_1}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_1}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11703977+sky130_fd_pr__nfet_01v8_lvt__voff_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.89325217+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_1}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_1}
+ etab = -0.0005
+ dsub = 0.40224308
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23453+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_1}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.011748
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00012443488
+ alpha1 = 0.0
+ beta0 = 21.191235
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26852+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_1}
+ kt2 = -0.037089
+ at = 49172.0
+ ute = -1.1197
+ ua1 = 2.0463e-9
+ ub1 = -1.8943e-18
+ uc1 = -9.1901e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.2 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 6.005e-06 wmin = 9.95e-07 wmax = 2.085e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.42802+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.53326
+ k2 = {-0.067164508+sky130_fd_pr__nfet_01v8_lvt__k2_diff_2}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {200550+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_2}
+ ua = {-9.7865e-010+sky130_fd_pr__nfet_01v8_lvt__ua_diff_2}
+ ub = {2.1353e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_2}
+ uc = 2.2350587e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_2}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.032501+sky130_fd_pr__nfet_01v8_lvt__u0_diff_2}
+ a0 = {1.9137+sky130_fd_pr__nfet_01v8_lvt__a0_diff_2}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.51517+sky130_fd_pr__nfet_01v8_lvt__ags_diff_2}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_2}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11023409+sky130_fd_pr__nfet_01v8_lvt__voff_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.8176398+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_2}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_2}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_2}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0075691
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.1734937e-5
+ alpha1 = 0.0
+ beta0 = 17.793363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25763+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_2}
+ kt2 = -0.036364
+ at = 58230.0
+ ute = -1.1808
+ ua1 = 1.9636e-9
+ ub1 = -1.466e-18
+ uc1 = 6.3418e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.3 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27009+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.6626
+ k2 = {-0.090794821+sky130_fd_pr__nfet_01v8_lvt__k2_diff_3}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {163560+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_3}
+ ua = {-2.1086e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_3}
+ ub = {2.2465e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_3}
+ uc = 9.6631013e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_3}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016895+sky130_fd_pr__nfet_01v8_lvt__u0_diff_3}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_3}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2458+sky130_fd_pr__nfet_01v8_lvt__ags_diff_3}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_3}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11291855+sky130_fd_pr__nfet_01v8_lvt__voff_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.7696915+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_3}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.048017216+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_3}
+ etab = -0.011685015
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33036+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_3}
+ pdiblc1 = 0.94998046
+ pdiblc2 = 0.0075387
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00018578676
+ alpha1 = 0.0
+ beta0 = 26.886024
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.29309+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_3}
+ kt2 = -0.0079249
+ at = 73790.0
+ ute = -1.6543
+ ua1 = -1.1099e-10
+ ub1 = 3.7483e-19
+ uc1 = -1.3108e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.4 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27187+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.73031
+ k2 = {-0.11367935+sky130_fd_pr__nfet_01v8_lvt__k2_diff_4}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {166950+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_4}
+ ua = {-2.2656e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_4}
+ ub = {2.4621e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_4}
+ uc = 3.0856067e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_4}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01582+sky130_fd_pr__nfet_01v8_lvt__u0_diff_4}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_4}
+ keta = {-0.10289323+sky130_fd_pr__nfet_01v8_lvt__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.0945+sky130_fd_pr__nfet_01v8_lvt__ags_diff_4}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_4}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.087984208+sky130_fd_pr__nfet_01v8_lvt__voff_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.5974262+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_4}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.074368062+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_4}
+ etab = -0.019985473
+ dsub = 0.33890038
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.24347+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_4}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.014403
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00047214078
+ alpha1 = 0.0
+ beta0 = 28.34264
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.30418+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_4}
+ kt2 = -0.020858
+ at = 74036.0
+ ute = -1.7595
+ ua1 = -2.3854e-10
+ ub1 = 4.4297e-19
+ uc1 = 1.0686e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.5 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.35153+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.60051
+ k2 = {-0.081814864+sky130_fd_pr__nfet_01v8_lvt__k2_diff_5}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {157610+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_5}
+ ua = {-2.1842e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_5}
+ ub = {2.5076e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_5}
+ uc = 4.1827914e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_5}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.018689+sky130_fd_pr__nfet_01v8_lvt__u0_diff_5}
+ a0 = {1.5147+sky130_fd_pr__nfet_01v8_lvt__a0_diff_5}
+ keta = {-0.027106406+sky130_fd_pr__nfet_01v8_lvt__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0+sky130_fd_pr__nfet_01v8_lvt__ags_diff_5}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_5}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11162446+sky130_fd_pr__nfet_01v8_lvt__voff_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.3345212+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_5}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0028690017+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_5}
+ etab = -0.0086070049
+ dsub = 0.34935946
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.55878+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_5}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.012315
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0014156647
+ alpha1 = 0.0
+ beta0 = 29.93198
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27123+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_5}
+ kt2 = -0.024486
+ at = 53140.0
+ ute = -1.0201
+ ua1 = 1.1382e-9
+ ub1 = -8.5913e-19
+ uc1 = 7.2256e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.6 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43518+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.47289
+ k2 = {-0.043650972+sky130_fd_pr__nfet_01v8_lvt__k2_diff_6}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {169100+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_6}
+ ua = {-1.841e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_6}
+ ub = {2.5267e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_6}
+ uc = 5.6759971e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_6}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.023061+sky130_fd_pr__nfet_01v8_lvt__u0_diff_6}
+ a0 = {0.97812+sky130_fd_pr__nfet_01v8_lvt__a0_diff_6}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.22649+sky130_fd_pr__nfet_01v8_lvt__ags_diff_6}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_6}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12282847+sky130_fd_pr__nfet_01v8_lvt__voff_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.0775821+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_6}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0027101593+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_6}
+ etab = -0.000125
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.32485+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_6}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0073456
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00014083814
+ alpha1 = 0.0
+ beta0 = 24.284439
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27068+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_6}
+ kt2 = -0.035797
+ at = 81396.0
+ ute = -1.1292
+ ua1 = 1.4609e-9
+ ub1 = -1.2921e-18
+ uc1 = -1.1706e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.7 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43687+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.43772
+ k2 = {-0.029563+sky130_fd_pr__nfet_01v8_lvt__k2_diff_7}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {78147+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_7}
+ ua = {-1.4872e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_7}
+ ub = {2.4924e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_7}
+ uc = 7.3523e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_7}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.027727+sky130_fd_pr__nfet_01v8_lvt__u0_diff_7}
+ a0 = {1.6103+sky130_fd_pr__nfet_01v8_lvt__a0_diff_7}
+ keta = {-0.18545+sky130_fd_pr__nfet_01v8_lvt__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {2.1454+sky130_fd_pr__nfet_01v8_lvt__ags_diff_7}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_7}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11610013+sky130_fd_pr__nfet_01v8_lvt__voff_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.99450786+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_7}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.00046581+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_7}
+ etab = -0.00047275
+ dsub = 0.78526904
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.09004+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_7}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.013228
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 4.7269108e-5
+ alpha1 = 0.0
+ beta0 = 20.812363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26519+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_7}
+ kt2 = -0.020948
+ at = 77133.0
+ ute = -1.1063
+ ua1 = 2.6996e-9
+ ub1 = -3.0597e-18
+ uc1 = -8.7824e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.8 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.44133+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.44248
+ k2 = {-0.023695+sky130_fd_pr__nfet_01v8_lvt__k2_diff_8}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {38113+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_8}
+ ua = {-1.2359e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_8}
+ ub = {2.4321e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_8}
+ uc = 8.8913e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_8}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.031741+sky130_fd_pr__nfet_01v8_lvt__u0_diff_8}
+ a0 = {1.8948+sky130_fd_pr__nfet_01v8_lvt__a0_diff_8}
+ keta = {-0.25181+sky130_fd_pr__nfet_01v8_lvt__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.8556+sky130_fd_pr__nfet_01v8_lvt__ags_diff_8}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_8}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11790286+sky130_fd_pr__nfet_01v8_lvt__voff_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.91173049+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_8}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_8}
+ etab = -0.00049217
+ dsub = 0.34422953
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.18376+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_8}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0079831
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00014201164
+ alpha1 = 0.0
+ beta0 = 21.469327
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25346+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_8}
+ kt2 = -0.036246
+ at = 42727.0
+ ute = -1.2103
+ ua1 = 2.2286e-9
+ ub1 = -2.4997e-18
+ uc1 = -5.3486e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.9 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 6.005e-06 wmin = 2.205e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43106+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.50407
+ k2 = {-0.055532161+sky130_fd_pr__nfet_01v8_lvt__k2_diff_9}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {169790+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_9}
+ ua = {-1.1001e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_9}
+ ub = {2.3643e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_9}
+ uc = 6.9010287e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_9}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.032806+sky130_fd_pr__nfet_01v8_lvt__u0_diff_9}
+ a0 = {1.6763+sky130_fd_pr__nfet_01v8_lvt__a0_diff_9}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.54695+sky130_fd_pr__nfet_01v8_lvt__ags_diff_9}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_9}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11480431+sky130_fd_pr__nfet_01v8_lvt__voff_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.82351304+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_9}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_9}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_9}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0067115
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.8823913e-5
+ alpha1 = 0.0
+ beta0 = 17.79575
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.2558+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_9}
+ kt2 = -0.03478
+ at = 318480.0
+ ute = -1.261
+ ua1 = 2.0849e-9
+ ub1 = -2.0887e-18
+ uc1 = -4.6822e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.10 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27581+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.64823
+ k2 = {-0.087406911+sky130_fd_pr__nfet_01v8_lvt__k2_diff_10}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {167000+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_10}
+ ua = {-2.3817e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_10}
+ ub = {2.6335e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_10}
+ uc = 2.7801766e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_10}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01552+sky130_fd_pr__nfet_01v8_lvt__u0_diff_10}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_10}
+ keta = {-0.17591628+sky130_fd_pr__nfet_01v8_lvt__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2474+sky130_fd_pr__nfet_01v8_lvt__ags_diff_10}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_10}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082362842+sky130_fd_pr__nfet_01v8_lvt__voff_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.1169257+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_10}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.079139243+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_10}
+ etab = 0.0
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16801+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_10}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.0058337
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00033433486
+ alpha1 = 0.0
+ beta0 = 27.963348
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.35576+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_10}
+ kt2 = -0.01165
+ at = 87087.0
+ ute = -1.6634
+ ua1 = 1.5299e-10
+ ub1 = -7.9485e-20
+ uc1 = -3.9208e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.11 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.28467+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.6924
+ k2 = {-0.10788872+sky130_fd_pr__nfet_01v8_lvt__k2_diff_11}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {163600+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_11}
+ ua = {-2.2472e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_11}
+ ub = {2.4923e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_11}
+ uc = 3.8992977e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_11}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.015982+sky130_fd_pr__nfet_01v8_lvt__u0_diff_11}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_11}
+ keta = {-0.11098086+sky130_fd_pr__nfet_01v8_lvt__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.1415+sky130_fd_pr__nfet_01v8_lvt__ags_diff_11}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_11}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.092416108+sky130_fd_pr__nfet_01v8_lvt__voff_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.6268174+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_11}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.080177319+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_11}
+ etab = -0.014812791
+ dsub = 0.33543563
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.21128+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_11}
+ pdiblc1 = 0.9970288
+ pdiblc2 = 0.012314
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00054476609
+ alpha1 = 0.0
+ beta0 = 28.649137
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.30247+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_11}
+ kt2 = -0.021837
+ at = 70444.0
+ ute = -1.7237
+ ua1 = -2.4904e-11
+ ub1 = 2.3083e-19
+ uc1 = -5.9776e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.12 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.35940117+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.59021354
+ k2 = {-0.083605504+sky130_fd_pr__nfet_01v8_lvt__k2_diff_12}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {161153.28+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_12}
+ ua = {-2.0759229e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_12}
+ ub = {2.4935708e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_12}
+ uc = 4.750487e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_12}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.020466323+sky130_fd_pr__nfet_01v8_lvt__u0_diff_12}
+ a0 = {1.4945377+sky130_fd_pr__nfet_01v8_lvt__a0_diff_12}
+ keta = {-0.033234596+sky130_fd_pr__nfet_01v8_lvt__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0+sky130_fd_pr__nfet_01v8_lvt__ags_diff_12}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_12}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11070501+sky130_fd_pr__nfet_01v8_lvt__voff_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.4204601+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_12}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0082066506+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_12}
+ etab = -0.018609296
+ dsub = 0.26417268
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.36231734+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_12}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.017097
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0020097469
+ alpha1 = 0.0
+ beta0 = 30.469968
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27101+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_12}
+ kt2 = -0.018574
+ at = 56390.0
+ ute = -1.6917
+ ua1 = 1.3075e-11
+ ub1 = 6.2584e-20
+ uc1 = -3.0151e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.13 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43296+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.43091
+ k2 = {-0.038466497+sky130_fd_pr__nfet_01v8_lvt__k2_diff_13}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {165480+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_13}
+ ua = {-1.2564e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_13}
+ ub = {2.0148e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_13}
+ uc = 4.8359e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_13}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.027923+sky130_fd_pr__nfet_01v8_lvt__u0_diff_13}
+ a0 = {1.8064+sky130_fd_pr__nfet_01v8_lvt__a0_diff_13}
+ keta = {-0.012102924+sky130_fd_pr__nfet_01v8_lvt__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.80816+sky130_fd_pr__nfet_01v8_lvt__ags_diff_13}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_13}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11113816+sky130_fd_pr__nfet_01v8_lvt__voff_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.235799+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_13}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {1e-5+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_13}
+ etab = -9.939227e-5
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.29415+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_13}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.010916
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00010964542
+ alpha1 = 0.0
+ beta0 = 23.745597
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25838+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_13}
+ kt2 = -0.024922
+ at = 71861.0
+ ute = -1.5423
+ ua1 = 2.9497e-10
+ ub1 = -6.6e-20
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.14 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.44085+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.43559
+ k2 = {-0.027932+sky130_fd_pr__nfet_01v8_lvt__k2_diff_14}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {73992+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_14}
+ ua = {-1.5313e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_14}
+ ub = {2.5578e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_14}
+ uc = 7.6172e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_14}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.028352+sky130_fd_pr__nfet_01v8_lvt__u0_diff_14}
+ a0 = {1.8312+sky130_fd_pr__nfet_01v8_lvt__a0_diff_14}
+ keta = {-0.16911+sky130_fd_pr__nfet_01v8_lvt__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {2.1115+sky130_fd_pr__nfet_01v8_lvt__ags_diff_14}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_14}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11555279+sky130_fd_pr__nfet_01v8_lvt__voff_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.0175057+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_14}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.00047259+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_14}
+ etab = -0.00047632
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.27339+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_14}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.012027
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.9804783e-5
+ alpha1 = 0.0
+ beta0 = 21.235324
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26442+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_14}
+ kt2 = -0.03563
+ at = 73755.0
+ ute = -1.1728
+ ua1 = 2.1764e-9
+ ub1 = -2.1594e-18
+ uc1 = -2.81e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.15 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.42701+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.49529
+ k2 = {-0.036322+sky130_fd_pr__nfet_01v8_lvt__k2_diff_15}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {48616+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_15}
+ ua = {-1.2502e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_15}
+ ub = {2.463e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_15}
+ uc = 9.6319e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_15}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.032149+sky130_fd_pr__nfet_01v8_lvt__u0_diff_15}
+ a0 = {1.9254+sky130_fd_pr__nfet_01v8_lvt__a0_diff_15}
+ keta = {-0.216+sky130_fd_pr__nfet_01v8_lvt__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.4285+sky130_fd_pr__nfet_01v8_lvt__ags_diff_15}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_15}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11135061+sky130_fd_pr__nfet_01v8_lvt__voff_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.91054759+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_15}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_15}
+ etab = -0.0005
+ dsub = 0.42135652
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.049306+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_15}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0087834
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00012909824
+ alpha1 = 0.0
+ beta0 = 21.317405
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.2646+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_15}
+ kt2 = -0.021848
+ at = 58230.0
+ ute = -1.2334
+ ua1 = 2.6296e-9
+ ub1 = -2.8755e-18
+ uc1 = -3.9499e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.16 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 6.005e-06 wmin = 3.665e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43669+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.40031
+ k2 = {-0.018155591+sky130_fd_pr__nfet_01v8_lvt__k2_diff_16}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {242950+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_16}
+ ua = {-1.2659e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_16}
+ ub = {2.5188e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_16}
+ uc = 7.0441e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_16}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.03202+sky130_fd_pr__nfet_01v8_lvt__u0_diff_16}
+ a0 = {1.917+sky130_fd_pr__nfet_01v8_lvt__a0_diff_16}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.59558+sky130_fd_pr__nfet_01v8_lvt__ags_diff_16}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_16}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11890341+sky130_fd_pr__nfet_01v8_lvt__voff_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.87044474+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_16}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_16}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.068446+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_16}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.006587
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 3.3789948e-5
+ alpha1 = 0.0
+ beta0 = 17.541356
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25403+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_16}
+ kt2 = -0.03469
+ at = 68095.0
+ ute = -1.1969
+ ua1 = 2.9253e-9
+ ub1 = -3.2731e-18
+ uc1 = -2.6978e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.17 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.265+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.68408
+ k2 = {-0.10092996+sky130_fd_pr__nfet_01v8_lvt__k2_diff_17}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159490+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_17}
+ ua = {-2.4839e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_17}
+ ub = {2.741e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_17}
+ uc = 2.0637e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_17}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0153+sky130_fd_pr__nfet_01v8_lvt__u0_diff_17}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_17}
+ keta = {-0.10107445+sky130_fd_pr__nfet_01v8_lvt__keta_diff_17}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2518+sky130_fd_pr__nfet_01v8_lvt__ags_diff_17}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_17}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11125373+sky130_fd_pr__nfet_01v8_lvt__voff_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.7361635+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_17}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.061320531+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_17}
+ etab = -0.011842783
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.26846+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_17}
+ pdiblc1 = 0.88733622
+ pdiblc2 = 0.00293
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00064658745
+ alpha1 = 0.0
+ beta0 = 29.169162
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27631+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_17}
+ kt2 = -0.011946
+ at = 74477.0
+ ute = -1.4241
+ ua1 = 5.2229e-10
+ ub1 = -4.6448e-19
+ uc1 = -2.5816e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.18 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.25199+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.70362
+ k2 = {-0.11306757+sky130_fd_pr__nfet_01v8_lvt__k2_diff_18}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {173730+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_18}
+ ua = {-2.4279e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_18}
+ ub = {2.6979e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_18}
+ uc = 3.5731e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_18}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.015453+sky130_fd_pr__nfet_01v8_lvt__u0_diff_18}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_18}
+ keta = {-0.084402688+sky130_fd_pr__nfet_01v8_lvt__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.1919+sky130_fd_pr__nfet_01v8_lvt__ags_diff_18}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_18}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.090318302+sky130_fd_pr__nfet_01v8_lvt__voff_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.7405461+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_18}
+ cit = 4.0851228e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.090968035+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_18}
+ etab = -0.016991172
+ dsub = 0.31798345
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.13722+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_18}
+ pdiblc1 = 0.99999854
+ pdiblc2 = 0.010137
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0014751785
+ alpha1 = 0.0
+ beta0 = 30.389816
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.30896+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_18}
+ kt2 = -0.031201
+ at = 83039.0
+ ute = -1.5889
+ ua1 = 2.8812e-10
+ ub1 = -1.6956e-19
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.19 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.36519+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.60123
+ k2 = {-0.086339858+sky130_fd_pr__nfet_01v8_lvt__k2_diff_19}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {163500+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_19}
+ ua = {-1.6939e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_19}
+ ub = {2.335e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_19}
+ uc = 6.2031292e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_19}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.026545+sky130_fd_pr__nfet_01v8_lvt__u0_diff_19}
+ a0 = {1.4463+sky130_fd_pr__nfet_01v8_lvt__a0_diff_19}
+ keta = {-0.035383769+sky130_fd_pr__nfet_01v8_lvt__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0+sky130_fd_pr__nfet_01v8_lvt__ags_diff_19}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_19}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11184994+sky130_fd_pr__nfet_01v8_lvt__voff_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.4864344+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_19}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0035852069+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_19}
+ etab = -0.056245935
+ dsub = 0.33950027
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.39248+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_19}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.014916
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0018437948
+ alpha1 = 0.0
+ beta0 = 30.497039
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24566+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_19}
+ kt2 = -0.025941
+ at = 48658.0
+ ute = -0.83944
+ ua1 = 2.537e-9
+ ub1 = -2.3672e-18
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.20 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43542+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.44399
+ k2 = {-0.036419634+sky130_fd_pr__nfet_01v8_lvt__k2_diff_20}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {181810+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_20}
+ ua = {-1.6157e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_20}
+ ub = {2.3385e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_20}
+ uc = 5.5832208e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_20}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.025086+sky130_fd_pr__nfet_01v8_lvt__u0_diff_20}
+ a0 = {1.5651+sky130_fd_pr__nfet_01v8_lvt__a0_diff_20}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.052001+sky130_fd_pr__nfet_01v8_lvt__ags_diff_20}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_20}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11448892+sky130_fd_pr__nfet_01v8_lvt__voff_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.2230329+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_20}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_20}
+ etab = -6.3091638e-5
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.38467+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_20}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0098886
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00011964049
+ alpha1 = 0.0
+ beta0 = 23.939816
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26556+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_20}
+ kt2 = -0.034425
+ at = 50265.0
+ ute = -1.0446
+ ua1 = 2.4044e-9
+ ub1 = -2.5541e-18
+ uc1 = -2.6056e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.21 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43416+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.4318
+ k2 = {-0.018853+sky130_fd_pr__nfet_01v8_lvt__k2_diff_21}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {72446+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_21}
+ ua = {-1.5035e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_21}
+ ub = {2.5663e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_21}
+ uc = 8.6552e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_21}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.028624+sky130_fd_pr__nfet_01v8_lvt__u0_diff_21}
+ a0 = {1.7527+sky130_fd_pr__nfet_01v8_lvt__a0_diff_21}
+ keta = {-0.22512+sky130_fd_pr__nfet_01v8_lvt__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {2.1654+sky130_fd_pr__nfet_01v8_lvt__ags_diff_21}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_21}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11469605+sky130_fd_pr__nfet_01v8_lvt__voff_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.0144745+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_21}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.00040654+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_21}
+ etab = -0.00045738
+ dsub = 0.62572026
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.23099+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_21}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.010409
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 6.3466057e-5
+ alpha1 = 0.0
+ beta0 = 21.398715
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25665+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_21}
+ kt2 = -0.012958
+ at = 72262.0
+ ute = -1.0102
+ ua1 = 3.2297e-9
+ ub1 = -3.6218e-18
+ uc1 = -8.1904e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.22 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43612+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.43039
+ k2 = {-0.02688+sky130_fd_pr__nfet_01v8_lvt__k2_diff_22}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {45491+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_22}
+ ua = {-1.2241e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_22}
+ ub = {2.5347e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_22}
+ uc = 7.2945e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_22}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.033495+sky130_fd_pr__nfet_01v8_lvt__u0_diff_22}
+ a0 = {1.996+sky130_fd_pr__nfet_01v8_lvt__a0_diff_22}
+ keta = {-0.18453+sky130_fd_pr__nfet_01v8_lvt__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.5415+sky130_fd_pr__nfet_01v8_lvt__ags_diff_22}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_22}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11589656+sky130_fd_pr__nfet_01v8_lvt__voff_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.8472686+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_22}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0005+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_22}
+ etab = -0.0005
+ dsub = 0.28297352
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2301+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_22}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0086915
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00012577963
+ alpha1 = 0.0
+ beta0 = 21.296605
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25363+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_22}
+ kt2 = -0.029655
+ at = 51378.0
+ ute = -1.1692
+ ua1 = 3.2521e-9
+ ub1 = -3.7668e-18
+ uc1 = -3.4748e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.23 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.42182+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.47213
+ k2 = {-0.040853+sky130_fd_pr__nfet_01v8_lvt__k2_diff_23}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {161140+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_23}
+ ua = {-1.2992e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_23}
+ ub = {2.474e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_23}
+ uc = 7.0152e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_23}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.03111+sky130_fd_pr__nfet_01v8_lvt__u0_diff_23}
+ a0 = {1.9564+sky130_fd_pr__nfet_01v8_lvt__a0_diff_23}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0.52266+sky130_fd_pr__nfet_01v8_lvt__ags_diff_23}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_23}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11559919+sky130_fd_pr__nfet_01v8_lvt__voff_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.7095479+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_23}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.08+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_23}
+ etab = -0.07
+ dsub = 0.56
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_23}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0047977
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.4345657e-5
+ alpha1 = 0.0
+ beta0 = 17.822982
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25364+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_23}
+ kt2 = -0.034423
+ at = 333080.0
+ ute = -1.0777
+ ua1 = 2.6823e-9
+ ub1 = -2.4433e-18
+ uc1 = -1.9223e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.24 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27938+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope2/sqrt(1))}
+ k1 = 0.62404
+ k2 = {-0.088152942+sky130_fd_pr__nfet_01v8_lvt__k2_diff_24}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {167110+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_24}
+ ua = {-2.1303e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_24}
+ ub = {2.5574e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_24}
+ uc = 6.7929e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_24}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.019161+sky130_fd_pr__nfet_01v8_lvt__u0_diff_24}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_24}
+ keta = {-0.18262975+sky130_fd_pr__nfet_01v8_lvt__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2511+sky130_fd_pr__nfet_01v8_lvt__ags_diff_24}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_24}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.077299489+sky130_fd_pr__nfet_01v8_lvt__voff_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.111486+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_24}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.079778236+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_24}
+ etab = 0.0
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16298+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_24}
+ pdiblc1 = 0.38459193
+ pdiblc2 = 0.0015537
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0003949429
+ alpha1 = 0.0
+ beta0 = 28.465005
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31794+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_24}
+ kt2 = -0.024372
+ at = 83749.0
+ ute = -1.6806
+ ua1 = 6.0118e-10
+ ub1 = -7.3201e-19
+ uc1 = 1.09e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.25 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.25974+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.69852
+ k2 = {-0.11267749+sky130_fd_pr__nfet_01v8_lvt__k2_diff_25}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {171590+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_25}
+ ua = {-2.3908e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_25}
+ ub = {2.727e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_25}
+ uc = 4.1338e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_25}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.016097+sky130_fd_pr__nfet_01v8_lvt__u0_diff_25}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_25}
+ keta = {-0.11730913+sky130_fd_pr__nfet_01v8_lvt__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2038+sky130_fd_pr__nfet_01v8_lvt__ags_diff_25}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_25}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.085388395+sky130_fd_pr__nfet_01v8_lvt__voff_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.7166939+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_25}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.077442702+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_25}
+ etab = -0.014827305
+ dsub = 0.32190545
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.14833+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_25}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.013708
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0006435735
+ alpha1 = 0.0
+ beta0 = 28.998989
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31355+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_25}
+ kt2 = -0.0156
+ at = 79939.0
+ ute = -1.9039
+ ua1 = 1.8262e-11
+ ub1 = -1.2097e-19
+ uc1 = 1.8835e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.26 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.36448+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.5799
+ k2 = {-0.081312236+sky130_fd_pr__nfet_01v8_lvt__k2_diff_26}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {164010+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_26}
+ ua = {-1.9394e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_26}
+ ub = {2.4942e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_26}
+ uc = 5.4304177e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_26}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.023448+sky130_fd_pr__nfet_01v8_lvt__u0_diff_26}
+ a0 = {1.6132+sky130_fd_pr__nfet_01v8_lvt__a0_diff_26}
+ keta = {-0.0046409768+sky130_fd_pr__nfet_01v8_lvt__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0+sky130_fd_pr__nfet_01v8_lvt__ags_diff_26}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_26}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.10972446+sky130_fd_pr__nfet_01v8_lvt__voff_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.4549256+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_26}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0057719981+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_26}
+ etab = -0.027300733
+ dsub = 0.27015818
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.38014+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_26}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.013941
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0028629629
+ alpha1 = 0.0
+ beta0 = 31.268363
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27285+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_26}
+ kt2 = -0.021644
+ at = 55216.0
+ ute = -1.6671
+ ua1 = 4.9023e-10
+ ub1 = -7.0183e-19
+ uc1 = -3.6538e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.27 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.43055+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.4297
+ k2 = {-0.031909522+sky130_fd_pr__nfet_01v8_lvt__k2_diff_27}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {131150+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_27}
+ ua = {-1.8013e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_27}
+ ub = {2.5802e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_27}
+ uc = 6.4626e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_27}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.024337+sky130_fd_pr__nfet_01v8_lvt__u0_diff_27}
+ a0 = {1.4583+sky130_fd_pr__nfet_01v8_lvt__a0_diff_27}
+ keta = {-0.0093611521+sky130_fd_pr__nfet_01v8_lvt__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.3295+sky130_fd_pr__nfet_01v8_lvt__ags_diff_27}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_27}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11440866+sky130_fd_pr__nfet_01v8_lvt__voff_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.1323146+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_27}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {1e-5+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_27}
+ etab = -6.2466101e-5
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.51701+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_27}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.01052
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00015972238
+ alpha1 = 0.0
+ beta0 = 24.379967
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26292+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_27}
+ kt2 = -0.025167
+ at = 72155.0
+ ute = -1.0156
+ ua1 = 2.3891e-9
+ ub1 = -2.5035e-18
+ uc1 = 8.5804e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.28 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.42624+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.47969
+ k2 = {-0.045764+sky130_fd_pr__nfet_01v8_lvt__k2_diff_28}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {91661+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_28}
+ ua = {-1.1877e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_28}
+ ub = {2.3166e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_28}
+ uc = 2.5191e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_28}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.032613+sky130_fd_pr__nfet_01v8_lvt__u0_diff_28}
+ a0 = {1.5598+sky130_fd_pr__nfet_01v8_lvt__a0_diff_28}
+ keta = {-0.13+sky130_fd_pr__nfet_01v8_lvt__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.7587+sky130_fd_pr__nfet_01v8_lvt__ags_diff_28}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_28}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.13015687+sky130_fd_pr__nfet_01v8_lvt__voff_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {0.81374728+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_28}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {6.4148e-005+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_28}
+ etab = 0.0
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.24428+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_28}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.011485
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 8.8408382e-5
+ alpha1 = 0.0
+ beta0 = 21.901006
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.25554+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_28}
+ kt2 = -0.031752
+ at = 85042.0
+ ute = -1.0564
+ ua1 = 2.108e-9
+ ub1 = -1.8965e-18
+ uc1 = 3.783e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.29 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.21757+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.7181
+ k2 = {-0.092615+sky130_fd_pr__nfet_01v8_lvt__k2_diff_29}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {155580+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_29}
+ ua = {-2.3305e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_29}
+ ub = {2.5738e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_29}
+ uc = 4.8634e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_29}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.014411+sky130_fd_pr__nfet_01v8_lvt__u0_diff_29}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_29}
+ keta = {-0.13135+sky130_fd_pr__nfet_01v8_lvt__keta_diff_29}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2431+sky130_fd_pr__nfet_01v8_lvt__ags_diff_29}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_29}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082600814+sky130_fd_pr__nfet_01v8_lvt__voff_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.908064+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_29}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.029174+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_29}
+ etab = -0.0020741
+ dsub = 0.26003878
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.36625+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_29}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.01172
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00012695724
+ alpha1 = 0.0
+ beta0 = 26.338346
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31729+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_29}
+ kt2 = -0.019491
+ at = 74483.0
+ ute = -1.724
+ ua1 = -2.2727e-10
+ ub1 = 3.4823e-19
+ uc1 = 1.9015e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.30 nmos
* DC IV MOS Parameters
+ lmin = 1.75e-07 lmax = 1.85e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.33106+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.69124
+ k2 = {-0.09867298+sky130_fd_pr__nfet_01v8_lvt__k2_diff_30}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {164730+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_30}
+ ua = {-1.7974e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_30}
+ ub = {2.1449e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_30}
+ uc = 6.5686e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_30}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.021618+sky130_fd_pr__nfet_01v8_lvt__u0_diff_30}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_30}
+ keta = {0+sky130_fd_pr__nfet_01v8_lvt__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.0994+sky130_fd_pr__nfet_01v8_lvt__ags_diff_30}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_30}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.12227844+sky130_fd_pr__nfet_01v8_lvt__voff_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.2673229+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_30}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.07268068+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_30}
+ etab = -0.031401879
+ dsub = 0.31809498
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.31119+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_30}
+ pdiblc1 = 0.039
+ pdiblc2 = 0.012343
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00050448511
+ alpha1 = 0.0
+ beta0 = 28.596405
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.26906+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_30}
+ kt2 = -0.029955
+ at = 69730.0
+ ute = -1.7417
+ ua1 = -8.226e-11
+ ub1 = 1.8785e-19
+ uc1 = -5.7596e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.31 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.45e-07 wmax = 5.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.21837+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.7181
+ k2 = {-0.092615+sky130_fd_pr__nfet_01v8_lvt__k2_diff_31}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {166030+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_31}
+ ua = {-2.2839e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_31}
+ ub = {2.8188e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_31}
+ uc = 2.8482e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_31}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.015105+sky130_fd_pr__nfet_01v8_lvt__u0_diff_31}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_31}
+ keta = {-0.063+sky130_fd_pr__nfet_01v8_lvt__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2431+sky130_fd_pr__nfet_01v8_lvt__ags_diff_31}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_31}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.0826+sky130_fd_pr__nfet_01v8_lvt__voff_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.908+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_31}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.029174+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_31}
+ etab = -0.0020741
+ dsub = 0.26003878
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.36625+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_31}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.01172
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 2.9e-6
+ alpha1 = 0.0
+ beta0 = 18.964
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31729+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_31}
+ kt2 = -0.019491
+ at = 84911.0
+ ute = -1.724
+ ua1 = -3.3636e-10
+ ub1 = 3.4823e-19
+ uc1 = 1.9015e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.32 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 6.35e-07 wmax = 6.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.22857+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.7181
+ k2 = {-0.092615+sky130_fd_pr__nfet_01v8_lvt__k2_diff_32}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {155580+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_32}
+ ua = {-2.3305e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_32}
+ ub = {2.5738e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_32}
+ uc = 4.8634e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_32}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.014411+sky130_fd_pr__nfet_01v8_lvt__u0_diff_32}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_32}
+ keta = {-0.063048+sky130_fd_pr__nfet_01v8_lvt__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2431+sky130_fd_pr__nfet_01v8_lvt__ags_diff_32}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_32}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082601+sky130_fd_pr__nfet_01v8_lvt__voff_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.9081+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_32}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.029174+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_32}
+ etab = -0.0020741
+ dsub = 0.26003878
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.31362+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_32}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.018049
+ pdiblcb = 0.0
+ drout = 1.0484
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 5.0783e-6
+ alpha1 = 0.0
+ beta0 = 20.017
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.33129+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_32}
+ kt2 = -0.019491
+ at = 82000.0
+ ute = -1.724
+ ua1 = -2.2727e-10
+ ub1 = 3.4823e-19
+ uc1 = 1.9015e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.33 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 8.35e-07 wmax = 8.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.22357+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.7181
+ k2 = {-0.092615+sky130_fd_pr__nfet_01v8_lvt__k2_diff_33}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159000+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33}
+ ua = {-2.3305e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_33}
+ ub = {2.6138e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_33}
+ uc = 4.8634e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.014411+sky130_fd_pr__nfet_01v8_lvt__u0_diff_33}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_33}
+ keta = {-0.10781+sky130_fd_pr__nfet_01v8_lvt__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2431+sky130_fd_pr__nfet_01v8_lvt__ags_diff_33}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_33}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082600814+sky130_fd_pr__nfet_01v8_lvt__voff_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.908064+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.029174+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33}
+ etab = -0.0020741
+ dsub = 0.26003878
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.018752
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.6174e-6
+ alpha1 = 0.0
+ beta0 = 20.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31729+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33}
+ kt2 = -0.019491
+ at = 77462.0
+ ute = -1.724
+ ua1 = -2.2727e-10
+ ub1 = 3.4823e-19
+ uc1 = 1.9015e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.34 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 1.645e-06 wmax = 1.655e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27581+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.64823
+ k2 = {-0.087406911+sky130_fd_pr__nfet_01v8_lvt__k2_diff_34}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {167000+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_34}
+ ua = {-2.3817e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_34}
+ ub = {2.6335e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_34}
+ uc = 2.7801766e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_34}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01552+sky130_fd_pr__nfet_01v8_lvt__u0_diff_34}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_34}
+ keta = {-0.17591628+sky130_fd_pr__nfet_01v8_lvt__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2474+sky130_fd_pr__nfet_01v8_lvt__ags_diff_34}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_34}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082362842+sky130_fd_pr__nfet_01v8_lvt__voff_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.1169257+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_34}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.079139243+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_34}
+ etab = 0.0
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16801+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_34}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.0058337
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00033433486
+ alpha1 = 0.0
+ beta0 = 27.963348
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.35576+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_34}
+ kt2 = -0.01165
+ at = 87087.0
+ ute = -1.6634
+ ua1 = 1.5299e-10
+ ub1 = -7.9485e-20
+ uc1 = -3.9208e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.35 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 3.005e-06 wmax = 3.015e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.27581+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.64823
+ k2 = {-0.087406911+sky130_fd_pr__nfet_01v8_lvt__k2_diff_35}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {167000+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_35}
+ ua = {-2.3817e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_35}
+ ub = {2.6335e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_35}
+ uc = 2.7801766e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_35}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.01552+sky130_fd_pr__nfet_01v8_lvt__u0_diff_35}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_35}
+ keta = {-0.17591628+sky130_fd_pr__nfet_01v8_lvt__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2474+sky130_fd_pr__nfet_01v8_lvt__ags_diff_35}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_35}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082362842+sky130_fd_pr__nfet_01v8_lvt__voff_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.1169257+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_35}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.079139243+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_35}
+ etab = 0.0
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.16801+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_35}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.0058337
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00033433486
+ alpha1 = 0.0
+ beta0 = 27.963348
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.35576+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_35}
+ kt2 = -0.01165
+ at = 87087.0
+ ute = -1.6634
+ ua1 = 1.5299e-10
+ ub1 = -7.9485e-20
+ uc1 = -3.9208e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.36 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.265+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.68408
+ k2 = {-0.10092996+sky130_fd_pr__nfet_01v8_lvt__k2_diff_36}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159490+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_36}
+ ua = {-2.4839e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_36}
+ ub = {2.741e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_36}
+ uc = 2.0637e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_36}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.0153+sky130_fd_pr__nfet_01v8_lvt__u0_diff_36}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_36}
+ keta = {-0.10107445+sky130_fd_pr__nfet_01v8_lvt__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2518+sky130_fd_pr__nfet_01v8_lvt__ags_diff_36}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_36}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11125373+sky130_fd_pr__nfet_01v8_lvt__voff_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.7361635+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_36}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.061320531+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_36}
+ etab = -0.011842783
+ dsub = 0.26
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.26846+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_36}
+ pdiblc1 = 0.88733622
+ pdiblc2 = 0.00293
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.00064658745
+ alpha1 = 0.0
+ beta0 = 29.169162
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.27631+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_36}
+ kt2 = -0.011946
+ at = 74477.0
+ ute = -1.4241
+ ua1 = 5.2229e-10
+ ub1 = -4.6448e-19
+ uc1 = -2.5816e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.37 nmos
* DC IV MOS Parameters
+ lmin = 2.45e-07 lmax = 2.55e-07 wmin = 5.045e-06 wmax = 5.055e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.36519+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.60123
+ k2 = {-0.086339858+sky130_fd_pr__nfet_01v8_lvt__k2_diff_37}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {163500+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_37}
+ ua = {-1.6939e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_37}
+ ub = {2.335e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_37}
+ uc = 6.2031292e-11
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_37}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.026545+sky130_fd_pr__nfet_01v8_lvt__u0_diff_37}
+ a0 = {1.4463+sky130_fd_pr__nfet_01v8_lvt__a0_diff_37}
+ keta = {-0.035383769+sky130_fd_pr__nfet_01v8_lvt__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {0+sky130_fd_pr__nfet_01v8_lvt__ags_diff_37}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_37}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.11184994+sky130_fd_pr__nfet_01v8_lvt__voff_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.4864344+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_37}
+ cit = 5.0e-6
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.0035852069+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_37}
+ etab = -0.056245935
+ dsub = 0.33950027
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.39248+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_37}
+ pdiblc1 = 0.39
+ pdiblc2 = 0.014916
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 0.0018437948
+ alpha1 = 0.0
+ beta0 = 30.497039
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.24566+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_37}
+ kt2 = -0.025941
+ at = 48658.0
+ ute = -0.83944
+ ua1 = 2.537e-9
+ ub1 = -2.3672e-18
+ uc1 = 0.0
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_01v8_lvt.38 nmos
* DC IV MOS Parameters
+ lmin = 1.45e-07 lmax = 1.55e-07 wmin = 7.35e-07 wmax = 7.45e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.148e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {1.2025e-008+sky130_fd_pr__nfet_01v8_lvt__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -1.33e-8
+ dwb = -1.08e-8
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = -3.0e-7
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 0.0
+ xn = 0.0
+ rnoia = 0.912
+ rnoib = 0.26
+ tnoia = 2.5e+7
+ tnoib = 9.9e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.148e-009*sky130_fd_pr__nfet_01v8_lvt__toxe_mult+MC_MM_SWITCH*(4.148e-09*sky130_fd_pr__nfet_01v8_lvt__toxe_mult*(sky130_fd_pr__nfet_01v8_lvt__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_01v8_lvt__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.22357+sky130_fd_pr__nfet_01v8_lvt__vth0_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__vth0_slope1/sqrt(1))}
+ k1 = 0.7181
+ k2 = {-0.092615+sky130_fd_pr__nfet_01v8_lvt__k2_diff_33}
+ k3 = 1.65
+ dvt0 = 0.07665
+ dvt1 = 0.1252
+ dvt2 = -0.05637
+ dvt0w = 0.0
+ dvt1w = 5300000.0
+ dvt2w = -0.032
+ w0 = 1.0e-7
+ k3b = 1.6
+ vfb = 0.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.3802e-7
+ lpeb = -4.9152e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {159000+sky130_fd_pr__nfet_01v8_lvt__vsat_diff_33}
+ ua = {-2.3305e-009+sky130_fd_pr__nfet_01v8_lvt__ua_diff_33}
+ ub = {2.6138e-018+sky130_fd_pr__nfet_01v8_lvt__ub_diff_33}
+ uc = 4.8634e-12
+ rdsw = {103.65+sky130_fd_pr__nfet_01v8_lvt__rdsw_diff_33}
+ prwb = 0.0
+ prwg = 0.0
+ wr = 1.0
+ u0 = {0.014411+sky130_fd_pr__nfet_01v8_lvt__u0_diff_33}
+ a0 = {0+sky130_fd_pr__nfet_01v8_lvt__a0_diff_33}
+ keta = {-0.10781+sky130_fd_pr__nfet_01v8_lvt__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.38689047
+ ags = {1.2431+sky130_fd_pr__nfet_01v8_lvt__ags_diff_33}
+ b0 = {0+sky130_fd_pr__nfet_01v8_lvt__b0_diff_33}
+ b1 = {0+sky130_fd_pr__nfet_01v8_lvt__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.082600814+sky130_fd_pr__nfet_01v8_lvt__voff_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {1.908064+sky130_fd_pr__nfet_01v8_lvt__nfactor_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_01v8_lvt__tvoff_diff_33}
+ cit = 1.0e-5
+ cdsc = 3.8556e-37
+ cdscb = -0.00011484
+ cdscd = 4.7984e-6
+ eta0 = {0.029174+sky130_fd_pr__nfet_01v8_lvt__eta0_diff_33}
+ etab = -0.0020741
+ dsub = 0.26003878
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33+sky130_fd_pr__nfet_01v8_lvt__pclm_diff_33}
+ pdiblc1 = 1.0
+ pdiblc2 = 0.018752
+ pdiblcb = 0.0
+ drout = 3.4946
+ pscbe1 = 4.5e+8
+ pscbe2 = 1.0e-8
+ pvag = 0.0
+ delta = 0.01
+ alpha0 = 7.6174e-6
+ alpha1 = 0.0
+ beta0 = 20.6
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = {1.4427e-015+sky130_fd_pr__nfet_01v8_lvt__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_01v8_lvt__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2.3e+9
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.148e-9
* Temperature Effects Parameters
+ kt1 = {-0.31729+sky130_fd_pr__nfet_01v8_lvt__kt1_diff_33}
+ kt2 = -0.019491
+ at = 77462.0
+ ute = -1.724
+ ua1 = -2.2727e-10
+ ub1 = 3.4823e-19
+ uc1 = 1.9015e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 9.0e+41
+ noib = 1.0e+27
+ noic = 800000000000.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 1.2
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.2928
+ jss = 0.0027500000000000003
+ jsws = 6.0e-10
+ xtis = 2.0
+ bvs = 11.9
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.0012287
+ tpbsw = 0.0
+ tpbswg = 0.0
+ tcj = 0.000792
+ tcjsw = 1.0e-5
+ tcjswg = 0.0
+ cgdo = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgso = {2.5889e-010*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgbo = 1.0e-14
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cgdl = {2.5e-011*sky130_fd_pr__nfet_01v8_lvt__overlap_mult}
+ cf = 1.0e-14
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {1.3469e-008+sky130_fd_pr__nfet_01v8_lvt__dlc_diff+sky130_fd_pr__nfet_01v8_lvt__dlc_rotweak}
+ dwc = {2.6e-008+sky130_fd_pr__nfet_01v8_lvt__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.38008
+ moin = 23.81
+ noff = 3.8661
+ voffcv = -0.16994
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.001209*sky130_fd_pr__nfet_01v8_lvt__ajunction_mult}
+ mjs = 0.42197
+ pbs = 0.7477
+ cjsws = {3.6224e-011*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjsws = 0.001
+ pbsws = 0.1
+ cjswgs = {2.0132e-010*sky130_fd_pr__nfet_01v8_lvt__pjunction_mult}
+ mjswgs = 0.8000
+ pbswgs = 0.79644
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ wlod = {0+sky130_fd_pr__nfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__nfet_01v8_lvt
