magic
tech gf180mcuC
timestamp 1661874280
<< nwell >>
rect 0 61 172 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 53 19 59 36
rect 85 19 91 36
rect 102 19 108 36
rect 124 19 130 36
rect 141 19 147 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 53 70 59 104
rect 85 70 91 104
rect 102 70 108 104
rect 124 70 130 104
rect 141 70 147 104
<< ndiff >>
rect 9 30 19 36
rect 9 21 11 30
rect 16 21 19 30
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 19 53 36
rect 59 34 69 36
rect 59 21 62 34
rect 67 21 69 34
rect 59 19 69 21
rect 75 27 85 36
rect 75 21 77 27
rect 82 21 85 27
rect 75 19 85 21
rect 91 34 102 36
rect 91 29 94 34
rect 99 29 102 34
rect 91 19 102 29
rect 108 27 124 36
rect 108 21 111 27
rect 116 21 124 27
rect 108 19 124 21
rect 130 34 141 36
rect 130 21 133 34
rect 138 21 141 34
rect 130 19 141 21
rect 147 34 162 36
rect 147 21 155 34
rect 160 21 162 34
rect 147 19 162 21
<< pdiff >>
rect 9 102 19 104
rect 9 77 11 102
rect 16 77 19 102
rect 9 70 19 77
rect 25 102 36 104
rect 25 72 28 102
rect 33 72 36 102
rect 25 70 36 72
rect 42 102 53 104
rect 42 72 45 102
rect 50 72 53 102
rect 42 70 53 72
rect 59 102 69 104
rect 59 72 62 102
rect 67 72 69 102
rect 59 70 69 72
rect 75 102 85 104
rect 75 72 77 102
rect 82 72 85 102
rect 75 70 85 72
rect 91 70 102 104
rect 108 102 124 104
rect 108 72 111 102
rect 121 72 124 102
rect 108 70 124 72
rect 130 102 141 104
rect 130 92 133 102
rect 138 92 141 102
rect 130 70 141 92
rect 147 102 162 104
rect 147 72 150 102
rect 160 72 162 102
rect 147 70 162 72
<< ndiffc >>
rect 11 21 16 30
rect 28 21 33 34
rect 62 21 67 34
rect 77 21 82 27
rect 94 29 99 34
rect 111 21 116 27
rect 133 21 138 34
rect 155 21 160 34
<< pdiffc >>
rect 11 77 16 102
rect 28 72 33 102
rect 45 72 50 102
rect 62 72 67 102
rect 77 72 82 102
rect 111 72 121 102
rect 133 92 138 102
rect 150 72 160 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 134 10 143 12
rect 134 5 136 10
rect 141 5 143 10
rect 134 3 143 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
rect 81 118 90 120
rect 81 113 83 118
rect 88 113 90 118
rect 81 111 90 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
rect 129 118 138 120
rect 129 113 131 118
rect 136 113 138 118
rect 129 111 138 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
rect 136 5 141 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
rect 107 113 112 118
rect 131 113 136 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 53 104 59 109
rect 85 104 91 109
rect 102 104 108 109
rect 124 104 130 109
rect 141 104 147 109
rect 19 67 25 70
rect 19 65 31 67
rect 19 59 23 65
rect 29 59 31 65
rect 19 57 31 59
rect 19 36 25 57
rect 36 52 42 70
rect 30 50 42 52
rect 53 51 59 70
rect 85 52 91 70
rect 30 44 32 50
rect 38 44 42 50
rect 30 42 42 44
rect 36 36 42 42
rect 47 49 59 51
rect 47 43 49 49
rect 55 43 59 49
rect 47 41 59 43
rect 78 50 91 52
rect 78 44 80 50
rect 86 44 91 50
rect 78 42 91 44
rect 53 36 59 41
rect 85 36 91 42
rect 102 48 108 70
rect 124 68 130 70
rect 124 66 136 68
rect 124 60 128 66
rect 134 60 136 66
rect 124 58 136 60
rect 102 46 112 48
rect 102 40 104 46
rect 110 40 112 46
rect 102 38 112 40
rect 102 36 108 38
rect 124 36 130 58
rect 141 52 147 70
rect 135 50 147 52
rect 135 44 137 50
rect 143 44 147 50
rect 135 42 147 44
rect 141 36 147 42
rect 19 14 25 19
rect 36 14 42 19
rect 53 14 59 19
rect 85 14 91 19
rect 102 14 108 19
rect 124 14 130 19
rect 141 14 147 19
<< polycontact >>
rect 23 59 29 65
rect 32 44 38 50
rect 49 43 55 49
rect 80 44 86 50
rect 128 60 134 66
rect 104 40 110 46
rect 137 44 143 50
<< metal1 >>
rect 0 118 172 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 131 118
rect 137 112 172 118
rect 0 111 172 112
rect 11 102 16 104
rect 11 76 16 77
rect 28 102 33 111
rect 8 70 10 76
rect 16 70 18 76
rect 28 70 33 72
rect 45 102 50 104
rect 11 30 16 70
rect 45 65 50 72
rect 62 102 67 111
rect 62 70 67 72
rect 77 102 82 111
rect 77 70 82 72
rect 111 102 121 104
rect 133 102 138 111
rect 133 90 138 92
rect 150 102 160 104
rect 111 70 121 72
rect 150 70 160 72
rect 21 59 23 65
rect 29 59 62 65
rect 68 59 70 65
rect 111 60 116 70
rect 126 60 128 66
rect 134 60 136 66
rect 155 64 160 70
rect 155 63 162 64
rect 30 44 32 50
rect 38 44 40 50
rect 47 43 49 49
rect 55 43 57 49
rect 49 37 55 43
rect 11 19 16 21
rect 28 34 33 36
rect 47 31 49 37
rect 55 31 57 37
rect 62 34 67 59
rect 94 55 121 60
rect 154 57 156 63
rect 162 57 164 63
rect 155 56 162 57
rect 78 44 80 50
rect 86 44 88 50
rect 28 12 33 21
rect 94 34 99 55
rect 115 50 135 55
rect 104 46 110 48
rect 130 44 137 50
rect 143 44 145 50
rect 104 38 110 40
rect 133 34 138 36
rect 62 19 67 21
rect 77 27 82 29
rect 94 27 99 29
rect 111 27 116 29
rect 82 21 111 22
rect 77 17 116 21
rect 133 12 138 21
rect 155 34 160 56
rect 155 19 160 21
rect 0 11 172 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 136 11
rect 142 5 172 11
rect 0 0 172 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 131 113 136 118
rect 136 113 137 118
rect 131 112 137 113
rect 10 70 16 76
rect 62 59 68 65
rect 128 60 134 66
rect 32 44 38 50
rect 49 31 55 37
rect 156 57 162 63
rect 80 44 86 50
rect 104 40 110 46
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 136 10 142 11
rect 136 5 141 10
rect 141 5 142 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 129 112 131 118
rect 137 112 139 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 8 76 18 77
rect 8 70 10 76
rect 16 70 18 76
rect 8 69 18 70
rect 126 66 136 67
rect 60 65 70 66
rect 126 65 128 66
rect 60 59 62 65
rect 68 60 128 65
rect 134 60 136 66
rect 68 59 136 60
rect 154 63 164 64
rect 60 58 70 59
rect 154 57 156 63
rect 162 57 164 63
rect 154 56 164 57
rect 30 50 40 51
rect 78 50 88 51
rect 30 44 32 50
rect 38 44 80 50
rect 86 44 88 50
rect 104 47 110 48
rect 30 43 40 44
rect 78 43 88 44
rect 103 46 111 47
rect 103 40 104 46
rect 110 40 111 46
rect 103 39 111 40
rect 48 37 56 38
rect 103 37 110 39
rect 47 31 49 37
rect 55 31 110 37
rect 48 30 56 31
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 135 11 143 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 134 5 136 11
rect 142 5 144 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 135 4 143 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 35 47 35 47 1 A
port 1 n
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 159 60 159 60 1 S
port 3 n
rlabel metal2 52 34 52 34 1 B
port 5 n
rlabel metal2 12 73 12 73 1 CO
port 4 n
<< end >>
