# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_xor2_1 0 0 ;
  SIZE 6.7 BY 6.15 ;
  SYMMETRY X Y ;
  SITE 9T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.1 2.2 1.6 2.5 ;
      LAYER MET2 ;
        RECT 1.1 2.2 1.6 2.5 ;
        RECT 1.15 2.15 1.55 2.55 ;
      LAYER VIA12 ;
        RECT 1.22 2.22 1.48 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.1 2.2 5.6 2.5 ;
        RECT 2.35 2 5.45 2.3 ;
      LAYER MET2 ;
        RECT 5.1 2.2 5.6 2.5 ;
        RECT 5.15 2.15 5.55 2.55 ;
      LAYER VIA12 ;
        RECT 5.22 2.22 5.48 2.48 ;
    END
  END B
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.7 0.6 ;
        RECT 5 0 5.25 1.75 ;
        RECT 1.4 0 1.65 1.8 ;
      LAYER MET2 ;
        RECT 5.25 0.25 5.75 0.55 ;
        RECT 5.3 0.2 5.7 0.6 ;
        RECT 4.05 0.25 4.55 0.55 ;
        RECT 4.1 0.2 4.5 0.6 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
        RECT 4.17 0.27 4.43 0.53 ;
        RECT 5.37 0.27 5.63 0.53 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 6.7 6.15 ;
        RECT 5 3.8 5.25 6.15 ;
        RECT 1.4 3.8 1.65 6.15 ;
      LAYER MET2 ;
        RECT 5.25 5.6 5.75 5.9 ;
        RECT 5.3 5.55 5.7 5.95 ;
        RECT 4.05 5.6 4.55 5.9 ;
        RECT 4.1 5.55 4.5 5.95 ;
        RECT 2.85 5.6 3.35 5.9 ;
        RECT 2.9 5.55 3.3 5.95 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
        RECT 2.97 5.62 3.23 5.88 ;
        RECT 4.17 5.62 4.43 5.88 ;
        RECT 5.37 5.62 5.63 5.88 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.05 1.4 3.55 1.7 ;
        RECT 3.15 1.3 3.45 1.75 ;
        RECT 3.2 0.95 3.45 1.75 ;
        RECT 3.05 4.15 3.55 4.45 ;
        RECT 3.2 4.15 3.45 5.2 ;
        RECT 3.15 4.15 3.45 4.55 ;
      LAYER MET2 ;
        RECT 3.05 1.35 3.55 1.75 ;
        RECT 3.1 4.1 3.5 4.5 ;
        RECT 3.15 1.35 3.45 4.55 ;
      LAYER VIA12 ;
        RECT 3.17 4.17 3.43 4.43 ;
        RECT 3.17 1.42 3.43 1.68 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.85 0.95 6.1 5.2 ;
      RECT 2.7 3.65 4.7 3.9 ;
      RECT 4.45 2.55 4.7 3.9 ;
      RECT 2.7 3.05 3 3.9 ;
      RECT 4.45 3.1 6.1 3.4 ;
      RECT 2.6 3.05 3.1 3.3 ;
      RECT 4.45 2.55 4.75 3.4 ;
      RECT 4.35 2.55 4.85 2.85 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 3.65 2.55 3.95 3.4 ;
      RECT 0.55 3 2.35 3.25 ;
      RECT 2.05 2.55 2.35 3.25 ;
      RECT 2.05 2.55 3.95 2.8 ;
  END
END gf180mcu_osu_sc_9T_xor2_1
