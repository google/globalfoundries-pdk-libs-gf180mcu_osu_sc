magic
tech gf180mcuC
timestamp 1659646792
<< nwell >>
rect 0 97 44 159
<< nmos >>
rect 19 16 25 33
<< pmos >>
rect 19 106 25 140
<< ndiff >>
rect 9 31 19 33
rect 9 18 11 31
rect 16 18 19 31
rect 9 16 19 18
rect 25 31 35 33
rect 25 18 28 31
rect 33 18 35 31
rect 25 16 35 18
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 35 140
rect 25 108 28 138
rect 33 108 35 138
rect 25 106 35 108
<< ndiffc >>
rect 11 18 16 31
rect 28 18 33 31
<< pdiffc >>
rect 11 108 16 138
rect 28 108 33 138
<< psubdiff >>
rect 9 7 18 9
rect 9 2 11 7
rect 16 2 18 7
rect 9 0 18 2
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
<< psubdiffcont >>
rect 11 2 16 7
<< nsubdiffcont >>
rect 11 149 16 154
<< polysilicon >>
rect 19 140 25 145
rect 19 48 25 106
rect 19 46 33 48
rect 19 41 26 46
rect 31 41 33 46
rect 19 39 33 41
rect 19 33 25 39
rect 19 11 25 16
<< polycontact >>
rect 26 41 31 46
<< metal1 >>
rect 0 154 44 159
rect 0 148 11 154
rect 17 148 44 154
rect 0 147 44 148
rect 11 138 16 147
rect 11 106 16 108
rect 28 138 33 140
rect 28 99 33 108
rect 26 93 28 99
rect 34 93 36 99
rect 28 92 33 93
rect 23 41 26 46
rect 31 41 33 46
rect 11 31 16 33
rect 11 9 16 18
rect 28 31 33 41
rect 28 16 33 18
rect 0 8 44 9
rect 0 2 11 8
rect 17 2 44 8
rect 0 -3 44 2
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 28 93 34 99
rect 11 7 17 8
rect 11 2 16 7
rect 16 2 17 7
<< metal2 >>
rect 10 154 18 155
rect 9 148 11 154
rect 17 148 19 154
rect 10 147 18 148
rect 26 99 36 100
rect 26 93 28 99
rect 34 93 36 99
rect 26 92 36 93
rect 10 8 18 9
rect 9 2 11 8
rect 17 2 19 8
rect 10 1 18 2
<< labels >>
rlabel metal2 14 5 14 5 1 GND
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 31 96 31 96 1 Y
port 2 n
<< end >>
