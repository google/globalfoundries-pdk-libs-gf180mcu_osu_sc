# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addh_1 0 0 ;
  SIZE 8.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 8.1 8.1 ;
        RECT 6.4 5.45 6.65 8.1 ;
        RECT 3.85 5.45 4.1 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.1 0.6 ;
        RECT 6.4 0 6.65 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 3.5 4.4 3.8 ;
        RECT 1.5 3.5 2 3.8 ;
      LAYER MET2 ;
        RECT 3.9 3.45 4.4 3.85 ;
        RECT 1.5 3.5 4.4 3.8 ;
        RECT 1.5 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.62 3.52 1.88 3.78 ;
        RECT 4.02 3.52 4.28 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 2.85 5.7 3.15 ;
        RECT 2.35 2.85 2.85 3.15 ;
      LAYER MET2 ;
        RECT 5.2 2.8 5.7 3.2 ;
        RECT 2.35 2.85 5.7 3.15 ;
        RECT 2.35 2.8 2.85 3.2 ;
      LAYER VIA12 ;
        RECT 2.47 2.87 2.73 3.13 ;
        RECT 5.32 2.87 5.58 3.13 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
        RECT 0.55 0.95 0.8 7.15 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.2 4.8 7.7 5.1 ;
        RECT 7.25 4.75 7.6 5.15 ;
        RECT 7.25 0.95 7.5 7.15 ;
      LAYER MET2 ;
        RECT 7.2 4.75 7.7 5.15 ;
      LAYER VIA12 ;
        RECT 7.32 4.82 7.58 5.08 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 6.05 4.75 6.55 5.15 ;
      RECT 3 4.75 3.5 5.15 ;
      RECT 3 4.8 6.55 5.1 ;
    LAYER VIA12 ;
      RECT 6.17 4.82 6.43 5.08 ;
      RECT 3.12 4.82 3.38 5.08 ;
    LAYER MET1 ;
      RECT 5.55 3.5 5.8 7.15 ;
      RECT 5.55 3.5 7 3.8 ;
      RECT 4.7 3.5 7 3.75 ;
      RECT 4.7 1.35 4.95 3.75 ;
      RECT 5.55 0.85 5.8 1.9 ;
      RECT 3.85 0.85 4.1 1.9 ;
      RECT 3.85 0.85 5.8 1.1 ;
      RECT 2.25 4.8 2.5 7.15 ;
      RECT 1.05 4.8 3.5 5.1 ;
      RECT 3.1 0.95 3.35 5.1 ;
      RECT 6.05 4.8 6.55 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addh_1
