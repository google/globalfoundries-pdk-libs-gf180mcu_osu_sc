VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addf_1 0 0 ;
  SIZE 14 BY 8.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 14 8.35 ;
        RECT 12.35 5.55 12.6 8.35 ;
        RECT 10.75 5.55 11 8.35 ;
        RECT 6.5 5.55 6.75 8.35 ;
        RECT 4.8 5.55 5.05 8.35 ;
        RECT 1.4 5.55 1.65 8.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14 0.7 ;
        RECT 12.35 0 12.6 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 6.5 0 6.75 1.55 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.7 3.6 9.2 3.9 ;
        RECT 4.6 3.6 5.1 3.9 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.6 9.2 3.9 ;
        RECT 8.75 3.55 9.15 3.95 ;
        RECT 4.65 3.55 5.05 3.95 ;
        RECT 0.65 3.55 1.05 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
        RECT 4.72 3.62 4.98 3.88 ;
        RECT 8.82 3.62 9.08 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.55 4.25 10.05 4.55 ;
        RECT 3.6 4.25 6.25 4.55 ;
        RECT 1.5 4.25 2 4.55 ;
      LAYER Metal2 ;
        RECT 5.75 4.25 10.05 4.55 ;
        RECT 9.6 4.2 10 4.6 ;
        RECT 5.8 4.2 6.2 4.6 ;
        RECT 1.5 4.25 4.1 4.55 ;
        RECT 3.65 4.2 4.05 4.6 ;
        RECT 1.55 4.2 1.95 4.6 ;
      LAYER Via1 ;
        RECT 1.62 4.27 1.88 4.53 ;
        RECT 3.72 4.27 3.98 4.53 ;
        RECT 5.87 4.27 6.13 4.53 ;
        RECT 9.67 4.27 9.93 4.53 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.05 2.3 10.55 2.6 ;
        RECT 6.65 2.3 7.15 2.6 ;
        RECT 2.35 2.95 2.85 3.25 ;
      LAYER Metal2 ;
        RECT 2.45 2.3 10.55 2.6 ;
        RECT 10.1 2.25 10.5 2.65 ;
        RECT 10.15 2.2 10.45 2.65 ;
        RECT 6.7 2.25 7.1 2.65 ;
        RECT 6.75 2.2 7.05 2.65 ;
        RECT 2.35 2.95 2.85 3.25 ;
        RECT 2.4 2.9 2.8 3.3 ;
        RECT 2.45 2.3 2.75 3.3 ;
      LAYER Via1 ;
        RECT 2.47 2.97 2.73 3.23 ;
        RECT 6.77 2.32 7.03 2.58 ;
        RECT 10.17 2.32 10.43 2.58 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.2 2.95 13.75 3.25 ;
        RECT 13.2 2.9 13.6 3.3 ;
        RECT 13.2 1.05 13.45 7.25 ;
      LAYER Metal2 ;
        RECT 13.25 2.95 13.75 3.25 ;
        RECT 13.3 2.9 13.7 3.3 ;
      LAYER Via1 ;
        RECT 13.37 2.97 13.63 3.23 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.6 4.25 12 4.55 ;
        RECT 11.6 1.05 11.85 7.25 ;
      LAYER Metal2 ;
        RECT 11.5 4.25 12 4.55 ;
        RECT 11.55 4.2 11.95 4.6 ;
      LAYER Via1 ;
        RECT 11.62 4.27 11.88 4.53 ;
    END
  END S
  OBS
    LAYER Metal2 ;
      RECT 12.5 2.9 12.9 3.3 ;
      RECT 7.5 2.9 7.9 3.3 ;
      RECT 7.45 2.95 12.95 3.25 ;
      RECT 12.55 2.85 12.85 3.3 ;
    LAYER Via1 ;
      RECT 12.57 2.97 12.83 3.23 ;
      RECT 7.57 2.97 7.83 3.23 ;
    LAYER Metal1 ;
      RECT 8.2 1.05 8.45 7.25 ;
      RECT 8.2 2.95 11.35 3.25 ;
      RECT 3.1 1.05 3.35 7.25 ;
      RECT 3.1 2.95 7.95 3.25 ;
      RECT 5.65 1.8 7.6 2.05 ;
      RECT 7.35 1.05 7.6 2.05 ;
      RECT 5.65 1.05 5.9 2.05 ;
      RECT 7.35 5.05 7.6 7.25 ;
      RECT 5.65 5.05 5.9 7.25 ;
      RECT 5.65 5.05 7.6 5.3 ;
      RECT 0.55 2.15 2.5 2.4 ;
      RECT 2.25 1.05 2.5 2.4 ;
      RECT 0.55 1.05 0.8 2.4 ;
      RECT 2.25 5.05 2.5 7.25 ;
      RECT 0.55 5.05 0.8 7.25 ;
      RECT 0.55 5.05 2.5 5.3 ;
      RECT 12.45 2.95 12.95 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addf_1

MACRO gf180mcu_osu_sc_gp12t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addh_1 0 0 ;
  SIZE 8.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 8.1 8.3 ;
        RECT 6.4 5.55 6.65 8.3 ;
        RECT 3.85 5.55 4.1 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 8.1 0.7 ;
        RECT 6.4 0 6.65 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.9 3.6 4.4 3.9 ;
        RECT 1.5 3.6 2 3.9 ;
      LAYER Metal2 ;
        RECT 3.9 3.55 4.4 3.95 ;
        RECT 1.5 3.6 4.4 3.9 ;
        RECT 1.5 3.55 2 3.95 ;
      LAYER Via1 ;
        RECT 1.62 3.62 1.88 3.88 ;
        RECT 4.02 3.62 4.28 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.2 2.95 5.7 3.25 ;
        RECT 2.35 2.95 2.85 3.25 ;
      LAYER Metal2 ;
        RECT 5.2 2.9 5.7 3.3 ;
        RECT 2.35 2.95 5.7 3.25 ;
        RECT 2.35 2.9 2.85 3.3 ;
      LAYER Via1 ;
        RECT 2.47 2.97 2.73 3.23 ;
        RECT 5.32 2.97 5.58 3.23 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 2.3 0.9 2.6 ;
        RECT 0.55 1.05 0.8 7.25 ;
      LAYER Metal2 ;
        RECT 0.4 2.25 0.9 2.65 ;
      LAYER Via1 ;
        RECT 0.52 2.32 0.78 2.58 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.2 4.9 7.7 5.2 ;
        RECT 7.25 4.85 7.6 5.25 ;
        RECT 7.25 1.05 7.5 7.25 ;
      LAYER Metal2 ;
        RECT 7.2 4.85 7.7 5.25 ;
      LAYER Via1 ;
        RECT 7.32 4.92 7.58 5.18 ;
    END
  END S
  OBS
    LAYER Metal2 ;
      RECT 6.05 4.85 6.55 5.25 ;
      RECT 3 4.85 3.5 5.25 ;
      RECT 3 4.9 6.55 5.2 ;
    LAYER Via1 ;
      RECT 6.17 4.92 6.43 5.18 ;
      RECT 3.12 4.92 3.38 5.18 ;
    LAYER Metal1 ;
      RECT 5.55 3.6 5.8 7.25 ;
      RECT 5.55 3.6 7 3.9 ;
      RECT 4.7 3.6 7 3.85 ;
      RECT 4.7 1.45 4.95 3.85 ;
      RECT 5.55 0.95 5.8 2 ;
      RECT 3.85 0.95 4.1 2 ;
      RECT 3.85 0.95 5.8 1.2 ;
      RECT 2.25 4.9 2.5 7.25 ;
      RECT 1.05 4.9 3.5 5.2 ;
      RECT 3.1 1.05 3.35 5.2 ;
      RECT 6.05 4.9 6.55 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addh_1

MACRO gf180mcu_osu_sc_gp12t3v3__and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__and2_1 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 2.1 0 2.5 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.55 1.1 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 2.95 2.4 3.25 ;
      LAYER Metal2 ;
        RECT 1.9 2.9 2.4 3.3 ;
      LAYER Via1 ;
        RECT 2.02 2.97 2.28 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 4.95 3.6 5.25 ;
        RECT 3.1 4.9 3.5 5.25 ;
        RECT 3.1 4.9 3.45 5.3 ;
        RECT 3.1 1.05 3.35 7.25 ;
      LAYER Metal2 ;
        RECT 3.1 4.9 3.6 5.3 ;
      LAYER Via1 ;
        RECT 3.22 4.97 3.48 5.23 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 2.35 4.2 2.85 4.6 ;
      RECT 1.3 4.2 1.8 4.6 ;
    LAYER Via1 ;
      RECT 2.47 4.27 2.73 4.53 ;
      RECT 1.42 4.27 1.68 4.53 ;
    LAYER Metal1 ;
      RECT 1.4 2 1.65 7.25 ;
      RECT 1.3 4.25 2.85 4.55 ;
      RECT 0.7 2 1.65 2.25 ;
      RECT 0.7 1.05 0.95 2.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__and2_1

MACRO gf180mcu_osu_sc_gp12t3v3__aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi21_1 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 1.4 6.3 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 2.95 0 3.2 1.9 ;
        RECT 0.7 0 0.95 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.55 1.1 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 4.25 2.1 4.55 ;
      LAYER Metal2 ;
        RECT 1.6 4.2 2.1 4.6 ;
      LAYER Via1 ;
        RECT 1.72 4.27 1.98 4.53 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.35 3.6 2.85 3.9 ;
      LAYER Metal2 ;
        RECT 2.35 3.55 2.85 3.95 ;
      LAYER Via1 ;
        RECT 2.47 3.62 2.73 3.88 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 4.9 3.5 5.2 ;
        RECT 3.1 2.65 3.35 7.25 ;
        RECT 2.1 2.65 3.35 2.9 ;
        RECT 2.1 1.05 2.35 2.9 ;
      LAYER Metal2 ;
        RECT 3 4.85 3.5 5.25 ;
      LAYER Via1 ;
        RECT 3.12 4.92 3.38 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 2.25 5.8 2.5 7.25 ;
      RECT 0.55 5.8 0.8 7.25 ;
      RECT 0.55 5.8 2.5 6.05 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi21_1

MACRO gf180mcu_osu_sc_gp12t3v3__aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi22_1 0 0 ;
  SIZE 5.35 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.35 8.3 ;
        RECT 1.4 6.3 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.35 0.7 ;
        RECT 3.5 0 3.75 1.9 ;
        RECT 0.7 0 0.95 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.55 1.1 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 4.25 2.1 4.55 ;
      LAYER Metal2 ;
        RECT 1.6 4.2 2.1 4.6 ;
      LAYER Via1 ;
        RECT 1.72 4.27 1.98 4.53 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.35 3.6 2.85 3.9 ;
      LAYER Metal2 ;
        RECT 2.35 3.55 2.85 3.95 ;
      LAYER Via1 ;
        RECT 2.47 3.62 2.73 3.88 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.3 4.25 3.8 4.55 ;
      LAYER Metal2 ;
        RECT 3.3 4.2 3.8 4.6 ;
      LAYER Via1 ;
        RECT 3.42 4.27 3.68 4.53 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.3 4.9 4.8 5.2 ;
        RECT 4.45 6.1 4.75 6.6 ;
        RECT 4.45 4.9 4.7 6.6 ;
        RECT 4.4 3.1 4.65 5.2 ;
        RECT 2.1 3.1 4.65 3.35 ;
        RECT 2.1 1.05 2.35 3.35 ;
        RECT 3 6.2 3.5 6.5 ;
        RECT 3.1 6.2 3.35 7.25 ;
      LAYER Metal2 ;
        RECT 4.35 6.15 4.85 6.55 ;
        RECT 3 6.2 4.85 6.5 ;
        RECT 3 6.15 3.5 6.55 ;
        RECT 4.3 4.85 4.8 5.25 ;
      LAYER Via1 ;
        RECT 3.12 6.22 3.38 6.48 ;
        RECT 4.42 4.92 4.68 5.18 ;
        RECT 4.47 6.22 4.73 6.48 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 3.95 5.7 4.2 7.25 ;
      RECT 2.25 5.7 2.5 7.25 ;
      RECT 0.55 5.7 0.8 7.25 ;
      RECT 0.55 5.7 4.2 5.95 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi22_1

MACRO gf180mcu_osu_sc_gp12t3v3__buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_1 0 0 ;
  SIZE 3.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.1 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.1 0.7 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.15 4.9 2.65 5.2 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.15 4.85 2.65 5.25 ;
      LAYER Via1 ;
        RECT 2.27 4.92 2.53 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_1

MACRO gf180mcu_osu_sc_gp12t3v3__buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_16 0 0 ;
  SIZE 15.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15.8 8.3 ;
        RECT 15 5.55 15.25 8.3 ;
        RECT 13.3 5.55 13.55 8.3 ;
        RECT 11.6 5.55 11.85 8.3 ;
        RECT 9.9 5.55 10.15 8.3 ;
        RECT 8.2 5.55 8.45 8.3 ;
        RECT 6.5 5.55 6.75 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15.8 0.7 ;
        RECT 15 0 15.25 1.9 ;
        RECT 13.3 0 13.55 1.9 ;
        RECT 11.6 0 11.85 1.9 ;
        RECT 9.9 0 10.15 1.9 ;
        RECT 8.2 0 8.45 1.9 ;
        RECT 6.5 0 6.75 1.9 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 14.05 4.9 14.55 5.2 ;
        RECT 14.15 1.05 14.4 7.25 ;
        RECT 2.25 4.95 14.4 5.25 ;
        RECT 2.25 2.15 14.4 2.4 ;
        RECT 12.45 1.05 12.7 7.25 ;
        RECT 10.75 1.05 11 7.25 ;
        RECT 9.05 1.05 9.3 7.25 ;
        RECT 7.35 1.05 7.6 7.25 ;
        RECT 5.65 1.05 5.9 7.25 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 14 4.95 14.55 5.25 ;
        RECT 14.05 4.85 14.55 5.25 ;
      LAYER Via1 ;
        RECT 14.17 4.92 14.43 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_16

MACRO gf180mcu_osu_sc_gp12t3v3__buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_2 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.15 4.9 2.65 5.2 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.15 4.85 2.65 5.25 ;
      LAYER Via1 ;
        RECT 2.27 4.92 2.53 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_2

MACRO gf180mcu_osu_sc_gp12t3v3__buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_4 0 0 ;
  SIZE 5.6 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.6 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.6 0.7 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.85 4.9 4.35 5.2 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 4.95 4.2 5.25 ;
        RECT 2.25 2.15 4.2 2.4 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 3.8 4.95 4.35 5.25 ;
        RECT 3.85 4.85 4.35 5.25 ;
      LAYER Via1 ;
        RECT 3.97 4.92 4.23 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_4

MACRO gf180mcu_osu_sc_gp12t3v3__buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__buf_8 0 0 ;
  SIZE 9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 9 8.3 ;
        RECT 8.2 5.55 8.45 8.3 ;
        RECT 6.5 5.55 6.75 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 9 0.7 ;
        RECT 8.2 0 8.45 1.9 ;
        RECT 6.5 0 6.75 1.9 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.25 4.9 7.75 5.2 ;
        RECT 7.35 1.05 7.6 7.25 ;
        RECT 2.25 4.95 7.6 5.25 ;
        RECT 2.25 2.15 7.6 2.4 ;
        RECT 5.65 1.05 5.9 7.25 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 7.2 4.95 7.75 5.25 ;
        RECT 7.25 4.85 7.75 5.25 ;
      LAYER Via1 ;
        RECT 7.37 4.92 7.63 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__buf_8

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_1 0 0 ;
  SIZE 3.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.1 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.1 0.7 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.15 4.9 2.65 5.2 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.15 4.85 2.65 5.25 ;
      LAYER Via1 ;
        RECT 2.27 4.92 2.53 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_1

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_16 0 0 ;
  SIZE 15.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15.8 8.3 ;
        RECT 15 5.55 15.25 8.3 ;
        RECT 13.3 5.55 13.55 8.3 ;
        RECT 11.6 5.55 11.85 8.3 ;
        RECT 9.9 5.55 10.15 8.3 ;
        RECT 8.2 5.55 8.45 8.3 ;
        RECT 6.5 5.55 6.75 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15.8 0.7 ;
        RECT 15 0 15.25 1.9 ;
        RECT 13.3 0 13.55 1.9 ;
        RECT 11.6 0 11.85 1.9 ;
        RECT 9.9 0 10.15 1.9 ;
        RECT 8.2 0 8.45 1.9 ;
        RECT 6.5 0 6.75 1.9 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 4.95 14.55 5.25 ;
        RECT 14.15 1.05 14.4 7.25 ;
        RECT 2.25 2.15 14.4 2.4 ;
        RECT 12.45 1.05 12.7 7.25 ;
        RECT 10.75 1.05 11 7.25 ;
        RECT 9.05 1.05 9.3 7.25 ;
        RECT 7.35 1.05 7.6 7.25 ;
        RECT 5.65 1.05 5.9 7.25 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 14.05 4.9 14.55 5.3 ;
        RECT 14 4.95 14.55 5.25 ;
      LAYER Via1 ;
        RECT 14.17 4.97 14.43 5.23 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_16

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_2 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.15 4.95 2.65 5.25 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.15 4.9 2.65 5.3 ;
      LAYER Via1 ;
        RECT 2.27 4.97 2.53 5.23 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_2

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_4 0 0 ;
  SIZE 5.6 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.6 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.6 0.7 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 4.95 4.35 5.25 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 2.15 4.2 2.4 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 3.85 4.9 4.35 5.3 ;
        RECT 3.8 4.95 4.35 5.25 ;
      LAYER Via1 ;
        RECT 3.97 4.97 4.23 5.23 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_4

MACRO gf180mcu_osu_sc_gp12t3v3__clkbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkbuf_8 0 0 ;
  SIZE 9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 9 8.3 ;
        RECT 8.2 5.55 8.45 8.3 ;
        RECT 6.5 5.55 6.75 8.3 ;
        RECT 4.8 5.55 5.05 8.3 ;
        RECT 3.1 5.55 3.35 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 9 0.7 ;
        RECT 8.2 0 8.45 1.9 ;
        RECT 6.5 0 6.75 1.9 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 4.95 7.75 5.25 ;
        RECT 7.35 1.05 7.6 7.25 ;
        RECT 2.25 2.15 7.6 2.4 ;
        RECT 5.65 1.05 5.9 7.25 ;
        RECT 3.95 1.05 4.2 7.25 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 7.25 4.9 7.75 5.3 ;
        RECT 7.2 4.95 7.75 5.25 ;
      LAYER Via1 ;
        RECT 7.37 4.97 7.63 5.23 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3 2 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__clkbuf_8

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_1 0 0 ;
  SIZE 2.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.2 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.2 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 3.6 1.8 3.9 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 1.3 3.55 1.8 3.95 ;
      LAYER Via1 ;
        RECT 1.42 3.62 1.68 3.88 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_1

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_16 0 0 ;
  SIZE 15 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15 8.3 ;
        RECT 14.15 5.55 14.4 8.3 ;
        RECT 12.45 5.55 12.7 8.3 ;
        RECT 10.75 5.55 11 8.3 ;
        RECT 9.05 5.55 9.3 8.3 ;
        RECT 7.35 5.55 7.6 8.3 ;
        RECT 5.65 5.55 5.9 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15 0.7 ;
        RECT 14.15 0 14.4 1.9 ;
        RECT 12.45 0 12.7 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 9.05 0 9.3 1.9 ;
        RECT 7.35 0 7.6 1.9 ;
        RECT 5.65 0 5.9 1.9 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.3 1.05 13.55 7.25 ;
        RECT 1.4 4.55 13.55 4.8 ;
        RECT 13.15 4.45 13.55 4.8 ;
        RECT 1.4 2.15 13.55 2.4 ;
        RECT 11.6 1.05 11.85 7.25 ;
        RECT 9.9 1.05 10.15 7.25 ;
        RECT 8.2 1.05 8.45 7.25 ;
        RECT 6.5 1.05 6.75 7.25 ;
        RECT 4.8 1.05 5.05 7.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 13.15 4.45 13.65 4.85 ;
      LAYER Via1 ;
        RECT 13.27 4.52 13.53 4.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_16

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_2 0 0 ;
  SIZE 3.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.2 8.3 ;
        RECT 2.3 5.55 2.55 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.2 0.7 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 3.6 1.15 3.9 ;
      LAYER Metal2 ;
        RECT 0.65 3.55 1.15 3.95 ;
      LAYER Via1 ;
        RECT 0.77 3.62 1.03 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.4 4.5 2 4.8 ;
        RECT 1.4 4.35 1.85 4.9 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 1.5 4.45 2 4.85 ;
      LAYER Via1 ;
        RECT 1.62 4.52 1.88 4.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_2

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_4 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 4.55 3.35 4.8 ;
        RECT 2.95 4.45 3.35 4.8 ;
        RECT 1.4 2.15 3.35 2.4 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 2.95 4.45 3.45 4.85 ;
      LAYER Via1 ;
        RECT 3.07 4.52 3.33 4.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_4

MACRO gf180mcu_osu_sc_gp12t3v3__clkinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__clkinv_8 0 0 ;
  SIZE 8.15 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 8.15 8.3 ;
        RECT 7.35 5.55 7.6 8.3 ;
        RECT 5.65 5.55 5.9 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 8.15 0.7 ;
        RECT 7.35 0 7.6 1.9 ;
        RECT 5.65 0 5.9 1.9 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.5 1.05 6.75 7.25 ;
        RECT 1.4 4.55 6.75 4.8 ;
        RECT 6.35 4.45 6.75 4.8 ;
        RECT 1.4 2.15 6.75 2.4 ;
        RECT 4.8 1.05 5.05 7.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 6.35 4.45 6.85 4.85 ;
      LAYER Via1 ;
        RECT 6.47 4.52 6.73 4.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__clkinv_8

MACRO gf180mcu_osu_sc_gp12t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dff_1 0 0 ;
  SIZE 13 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 13 8.3 ;
        RECT 11.3 5.55 11.55 8.3 ;
        RECT 8.85 5.55 9.1 8.3 ;
        RECT 7.25 6.3 7.5 8.3 ;
        RECT 4.45 5.55 4.7 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 13 0.7 ;
        RECT 11.3 0 11.55 1.9 ;
        RECT 8.85 0 9.1 1.55 ;
        RECT 7.25 0 7.5 1.9 ;
        RECT 4.45 0 4.7 1.5 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 7.65 4.25 8.15 4.55 ;
        RECT 5.5 4.25 6.55 4.55 ;
        RECT 5.4 2.25 5.9 2.55 ;
        RECT 5.5 2.25 5.8 4.55 ;
        RECT 2.6 4.25 3.75 4.55 ;
        RECT 3.25 2.3 3.75 2.6 ;
        RECT 3.35 2.3 3.65 4.55 ;
      LAYER Metal2 ;
        RECT 3.25 4.25 8.15 4.55 ;
        RECT 7.7 4.2 8.1 4.6 ;
        RECT 6.05 4.2 6.55 4.6 ;
        RECT 3.25 4.2 3.7 4.6 ;
      LAYER Via1 ;
        RECT 3.37 4.27 3.63 4.53 ;
        RECT 6.17 4.27 6.43 4.53 ;
        RECT 7.77 4.27 8.03 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 3.6 2.4 3.9 ;
      LAYER Metal2 ;
        RECT 1.75 3.6 2.55 3.9 ;
        RECT 1.9 3.55 2.4 3.95 ;
      LAYER Via1 ;
        RECT 2.02 3.62 2.28 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12.15 4.9 12.65 5.25 ;
        RECT 12.15 4.85 12.6 5.25 ;
        RECT 12.15 1.05 12.4 7.25 ;
      LAYER Metal2 ;
        RECT 12.15 4.9 12.65 5.2 ;
        RECT 12.2 4.85 12.6 5.25 ;
      LAYER Via1 ;
        RECT 12.27 4.92 12.53 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.45 4.25 11.9 4.55 ;
        RECT 11.55 2.15 11.8 4.55 ;
        RECT 10.45 2.15 11.8 2.4 ;
        RECT 10.45 4.25 10.7 7.25 ;
        RECT 10.45 1.05 10.7 2.4 ;
      LAYER Metal2 ;
        RECT 11.4 4.25 11.9 4.55 ;
        RECT 11.45 4.2 11.85 4.6 ;
      LAYER Via1 ;
        RECT 11.52 4.27 11.78 4.53 ;
    END
  END QN
  OBS
    LAYER Metal2 ;
      RECT 6.75 4.85 7.15 5.25 ;
      RECT 6.7 4.9 9.9 5.2 ;
      RECT 9.6 2.95 9.9 5.2 ;
      RECT 10.7 2.9 11.1 3.3 ;
      RECT 9.6 2.95 11.15 3.25 ;
      RECT 9 1.75 9.4 2.15 ;
      RECT 8.5 1.8 9.45 2.1 ;
      RECT 5.8 1.6 6.2 2 ;
      RECT 5.75 1.65 8.8 1.95 ;
      RECT 5.75 1.75 9.4 1.95 ;
      RECT 8.05 2.9 8.45 3.3 ;
      RECT 6.1 2.9 6.5 3.3 ;
      RECT 6.05 2.95 8.55 3.25 ;
      RECT 6.8 3.55 7.2 3.95 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 4.1 2.25 4.5 2.65 ;
      RECT 0.45 2.25 0.85 2.65 ;
      RECT 0.4 2.3 4.55 2.6 ;
    LAYER Via1 ;
      RECT 10.77 2.97 11.03 3.23 ;
      RECT 9.07 1.82 9.33 2.08 ;
      RECT 8.12 2.97 8.38 3.23 ;
      RECT 6.87 3.62 7.13 3.88 ;
      RECT 6.82 4.92 7.08 5.18 ;
      RECT 6.17 2.97 6.43 3.23 ;
      RECT 5.87 1.67 6.13 1.93 ;
      RECT 4.17 2.32 4.43 2.58 ;
      RECT 0.52 2.32 0.78 2.58 ;
    LAYER Metal1 ;
      RECT 9.7 1.05 9.95 7.25 ;
      RECT 9.7 2.95 11.15 3.25 ;
      RECT 9.05 1.8 9.35 3.35 ;
      RECT 8.95 2.95 9.45 3.25 ;
      RECT 8.95 1.8 9.45 2.1 ;
      RECT 8.1 4.85 8.35 7.25 ;
      RECT 8.1 4.85 8.9 5.1 ;
      RECT 8.6 3.65 8.9 5.1 ;
      RECT 8.1 3.65 8.9 3.9 ;
      RECT 8.1 2.85 8.4 3.9 ;
      RECT 8.1 1.05 8.35 3.9 ;
      RECT 6.7 4.9 7.2 5.2 ;
      RECT 6.8 3.55 7.1 5.2 ;
      RECT 6.75 3.6 7.3 3.9 ;
      RECT 6.8 3.55 7.2 3.9 ;
      RECT 5.85 6.05 6.1 7.25 ;
      RECT 4.95 6.05 6.1 6.3 ;
      RECT 4.95 3.55 5.2 6.3 ;
      RECT 4.9 1.7 5.15 3.8 ;
      RECT 4.9 1.7 6.25 1.95 ;
      RECT 5.85 1.65 6.25 1.95 ;
      RECT 5.85 1.05 6.1 1.95 ;
      RECT 4.05 4.9 4.55 5.2 ;
      RECT 4.15 2.3 4.45 5.2 ;
      RECT 4.05 2.3 4.55 2.6 ;
      RECT 3.05 5.05 3.3 7.25 ;
      RECT 1.4 5.05 3.3 5.3 ;
      RECT 1.4 2.35 1.65 5.3 ;
      RECT 1.05 4.25 1.65 4.55 ;
      RECT 1.4 2.35 2.4 2.6 ;
      RECT 2 1.65 2.4 2.6 ;
      RECT 2 1.65 3.3 1.9 ;
      RECT 3.05 1.05 3.3 1.9 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.5 2.2 0.8 2.7 ;
      RECT 6.05 2.95 6.55 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dff_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffn_1 0 0 ;
  SIZE 14.25 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 14.25 8.3 ;
        RECT 12.55 5.55 12.8 8.3 ;
        RECT 9.95 5.55 10.35 8.3 ;
        RECT 7.25 6.3 7.5 8.3 ;
        RECT 4.45 5.55 4.7 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14.25 0.7 ;
        RECT 12.55 0 12.8 1.9 ;
        RECT 9.95 0 10.35 1.55 ;
        RECT 7.25 0 7.5 1.9 ;
        RECT 4.45 0 4.7 1.5 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 9.5 2.95 10 3.25 ;
        RECT 9.6 2.85 9.9 3.35 ;
      LAYER Metal2 ;
        RECT 9.5 2.95 10 3.25 ;
        RECT 9.55 2.9 9.95 3.3 ;
      LAYER Via1 ;
        RECT 9.62 2.97 9.88 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 3.6 2.4 3.9 ;
      LAYER Metal2 ;
        RECT 1.75 3.6 2.55 3.9 ;
        RECT 1.9 3.55 2.4 3.95 ;
      LAYER Via1 ;
        RECT 2.02 3.62 2.28 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.4 4.9 13.9 5.25 ;
        RECT 13.4 4.85 13.85 5.25 ;
        RECT 13.4 1.05 13.65 7.25 ;
      LAYER Metal2 ;
        RECT 13.4 4.9 13.9 5.2 ;
        RECT 13.45 4.85 13.85 5.25 ;
      LAYER Via1 ;
        RECT 13.52 4.92 13.78 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.7 4.25 13.15 4.55 ;
        RECT 12.8 2.15 13.05 4.55 ;
        RECT 11.7 2.15 13.05 2.4 ;
        RECT 11.7 4.25 11.95 7.25 ;
        RECT 11.7 1.05 11.95 2.4 ;
      LAYER Metal2 ;
        RECT 12.65 4.25 13.15 4.55 ;
        RECT 12.7 4.2 13.1 4.6 ;
      LAYER Via1 ;
        RECT 12.77 4.27 13.03 4.53 ;
    END
  END QN
  OBS
    LAYER Metal2 ;
      RECT 6.75 4.85 7.15 5.25 ;
      RECT 6.7 4.9 11.15 5.2 ;
      RECT 10.85 2.95 11.15 5.2 ;
      RECT 11.95 2.9 12.35 3.3 ;
      RECT 10.85 2.95 12.4 3.25 ;
      RECT 10.25 1.75 10.65 2.15 ;
      RECT 9.5 1.8 10.7 2.1 ;
      RECT 5.8 1.6 6.2 2 ;
      RECT 5.75 1.65 9.9 1.95 ;
      RECT 5.75 1.75 10.65 1.95 ;
      RECT 8.9 4.2 9.3 4.6 ;
      RECT 7.7 4.2 8.1 4.6 ;
      RECT 6.05 4.2 6.55 4.6 ;
      RECT 3.25 4.2 3.7 4.6 ;
      RECT 3.25 4.25 9.35 4.55 ;
      RECT 8.05 2.9 8.45 3.3 ;
      RECT 6.1 2.9 6.5 3.3 ;
      RECT 6.05 2.95 8.55 3.25 ;
      RECT 6.8 3.55 7.2 3.95 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 4.1 2.25 4.5 2.65 ;
      RECT 0.45 2.25 0.85 2.65 ;
      RECT 0.4 2.3 4.55 2.6 ;
    LAYER Via1 ;
      RECT 12.02 2.97 12.28 3.23 ;
      RECT 10.32 1.82 10.58 2.08 ;
      RECT 8.97 4.27 9.23 4.53 ;
      RECT 8.12 2.97 8.38 3.23 ;
      RECT 7.77 4.27 8.03 4.53 ;
      RECT 6.87 3.62 7.13 3.88 ;
      RECT 6.82 4.92 7.08 5.18 ;
      RECT 6.17 2.97 6.43 3.23 ;
      RECT 6.17 4.27 6.43 4.53 ;
      RECT 5.87 1.67 6.13 1.93 ;
      RECT 4.17 2.32 4.43 2.58 ;
      RECT 3.37 4.27 3.63 4.53 ;
      RECT 0.52 2.32 0.78 2.58 ;
    LAYER Metal1 ;
      RECT 10.95 1.05 11.2 7.25 ;
      RECT 10.95 2.95 12.4 3.25 ;
      RECT 10.3 1.8 10.6 5.3 ;
      RECT 10.2 4.9 10.7 5.2 ;
      RECT 10.2 1.8 10.7 2.1 ;
      RECT 9.1 5.55 9.35 7.25 ;
      RECT 8.95 1.7 9.25 5.8 ;
      RECT 9.1 1.05 9.35 1.95 ;
      RECT 8.1 4.85 8.35 7.25 ;
      RECT 8.1 4.85 8.7 5.1 ;
      RECT 8.4 3.65 8.7 5.1 ;
      RECT 8.1 2.85 8.4 3.9 ;
      RECT 8.1 1.05 8.35 3.9 ;
      RECT 6.7 4.9 7.2 5.2 ;
      RECT 6.8 3.6 7.1 5.2 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 5.5 4.25 6.55 4.55 ;
      RECT 5.5 2.25 5.8 4.55 ;
      RECT 5.4 2.25 5.9 2.55 ;
      RECT 5.85 6.05 6.1 7.25 ;
      RECT 4.95 6.05 6.1 6.3 ;
      RECT 4.95 3.55 5.2 6.3 ;
      RECT 4.9 1.7 5.15 3.8 ;
      RECT 4.9 1.7 6.25 1.95 ;
      RECT 5.85 1.65 6.25 1.95 ;
      RECT 5.85 1.05 6.1 1.95 ;
      RECT 4.05 4.9 4.55 5.2 ;
      RECT 4.15 2.3 4.45 5.2 ;
      RECT 4.05 2.3 4.55 2.6 ;
      RECT 2.6 4.25 3.75 4.55 ;
      RECT 3.35 2.3 3.65 4.55 ;
      RECT 3.25 2.3 3.75 2.6 ;
      RECT 3.05 5.05 3.3 7.25 ;
      RECT 1.4 5.05 3.3 5.3 ;
      RECT 1.4 2.35 1.65 5.3 ;
      RECT 1.05 4.25 1.65 4.55 ;
      RECT 1.4 2.35 2.4 2.6 ;
      RECT 2 1.65 2.4 2.6 ;
      RECT 2 1.65 3.3 1.9 ;
      RECT 3.05 1.05 3.3 1.9 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.5 2.2 0.8 2.7 ;
      RECT 7.65 4.25 8.15 4.55 ;
      RECT 6.05 2.95 6.55 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffr_1 0 0 ;
  SIZE 17.6 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 17.6 8.3 ;
        RECT 15.95 5.55 16.2 8.3 ;
        RECT 12.95 5.55 13.2 8.3 ;
        RECT 10.75 6.3 11 8.3 ;
        RECT 7.95 5.55 8.2 8.3 ;
        RECT 4.9 5.55 5.15 8.3 ;
        RECT 3.55 5.55 3.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 17.6 0.7 ;
        RECT 15.95 0 16.2 1.9 ;
        RECT 14.2 0 14.45 1.9 ;
        RECT 12.5 0 12.75 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 7.95 0 8.2 1.5 ;
        RECT 4.9 0 5.15 1.9 ;
        RECT 4 0 4.25 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 11.15 4.25 11.65 4.55 ;
        RECT 9 4.25 10.05 4.55 ;
        RECT 8.9 2.25 9.4 2.55 ;
        RECT 9 2.25 9.3 4.55 ;
        RECT 6.1 4.25 7.25 4.55 ;
        RECT 6.75 2.3 7.25 2.6 ;
        RECT 6.85 2.3 7.15 4.55 ;
      LAYER Metal2 ;
        RECT 6.75 4.25 11.65 4.55 ;
        RECT 11.2 4.2 11.6 4.6 ;
        RECT 9.55 4.2 10.05 4.6 ;
        RECT 6.75 4.2 7.2 4.6 ;
      LAYER Via1 ;
        RECT 6.87 4.27 7.13 4.53 ;
        RECT 9.67 4.27 9.93 4.53 ;
        RECT 11.27 4.27 11.53 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.4 3.6 5.9 3.9 ;
      LAYER Metal2 ;
        RECT 5.4 3.55 5.9 3.95 ;
      LAYER Via1 ;
        RECT 5.52 3.62 5.78 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.8 4.9 17.3 5.25 ;
        RECT 16.8 4.85 17.25 5.25 ;
        RECT 16.8 1.05 17.05 7.25 ;
      LAYER Metal2 ;
        RECT 16.8 4.9 17.3 5.2 ;
        RECT 16.85 4.85 17.25 5.25 ;
      LAYER Via1 ;
        RECT 16.92 4.92 17.18 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15.1 4.25 16.55 4.55 ;
        RECT 16.2 2.15 16.45 4.55 ;
        RECT 15.1 2.15 16.45 2.4 ;
        RECT 15.1 4.25 15.35 7.25 ;
        RECT 15.1 1.05 15.35 2.4 ;
      LAYER Metal2 ;
        RECT 16.05 4.25 16.55 4.55 ;
        RECT 16.1 4.2 16.5 4.6 ;
      LAYER Via1 ;
        RECT 16.17 4.27 16.43 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  OBS
    LAYER Metal2 ;
      RECT 15.35 2.9 15.75 3.3 ;
      RECT 15 2.95 15.8 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 13.75 2.2 14.35 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 13.75 1 14.05 2.6 ;
      RECT 2.75 1 14.05 1.3 ;
      RECT 12.4 2.2 12.9 2.6 ;
      RECT 12.4 1.65 12.8 2.6 ;
      RECT 9.3 1.6 9.7 2 ;
      RECT 9.25 1.65 12.8 1.95 ;
      RECT 12.45 4.85 12.85 5.25 ;
      RECT 10.25 4.85 10.65 5.25 ;
      RECT 10.2 4.9 12.9 5.2 ;
      RECT 11.55 2.9 11.95 3.3 ;
      RECT 9.6 2.9 10 3.3 ;
      RECT 9.55 2.95 12.05 3.25 ;
      RECT 10.3 3.55 10.7 3.95 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 7.6 2.25 8 2.65 ;
      RECT 3.85 2.25 4.35 2.65 ;
      RECT 3.85 2.3 8.05 2.6 ;
      RECT 14.25 4.85 14.75 5.25 ;
    LAYER Via1 ;
      RECT 15.42 2.97 15.68 3.23 ;
      RECT 14.37 4.92 14.63 5.18 ;
      RECT 13.97 2.27 14.23 2.53 ;
      RECT 12.52 2.27 12.78 2.53 ;
      RECT 12.52 4.92 12.78 5.18 ;
      RECT 11.62 2.97 11.88 3.23 ;
      RECT 10.37 3.62 10.63 3.88 ;
      RECT 10.32 4.92 10.58 5.18 ;
      RECT 9.67 2.97 9.93 3.23 ;
      RECT 9.37 1.67 9.63 1.93 ;
      RECT 7.67 2.32 7.93 2.58 ;
      RECT 3.97 2.32 4.23 2.58 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 14.35 2.95 14.6 7.25 ;
      RECT 12.5 4.8 12.8 5.3 ;
      RECT 12.5 4.9 14.75 5.2 ;
      RECT 13.35 2.95 15.8 3.25 ;
      RECT 13.35 1.05 13.6 3.25 ;
      RECT 11.6 4.85 11.85 7.25 ;
      RECT 11.6 4.85 12.15 5.1 ;
      RECT 11.9 3.65 12.15 5.1 ;
      RECT 11.6 2.85 11.9 3.9 ;
      RECT 11.6 1.05 11.85 3.9 ;
      RECT 10.2 4.9 10.7 5.2 ;
      RECT 10.3 3.6 10.6 5.2 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 9.35 6.05 9.6 7.25 ;
      RECT 8.45 6.05 9.6 6.3 ;
      RECT 8.45 3.55 8.7 6.3 ;
      RECT 8.4 1.7 8.65 3.8 ;
      RECT 8.4 1.7 9.75 1.95 ;
      RECT 9.35 1.65 9.75 1.95 ;
      RECT 9.35 1.05 9.6 1.95 ;
      RECT 7.55 4.9 8.05 5.2 ;
      RECT 7.65 2.3 7.95 5.2 ;
      RECT 7.55 2.3 8.05 2.6 ;
      RECT 6.55 5.05 6.8 7.25 ;
      RECT 4.9 5.05 6.8 5.3 ;
      RECT 4.9 2.35 5.15 5.3 ;
      RECT 3.85 4.25 5.15 4.55 ;
      RECT 4.9 2.35 5.9 2.6 ;
      RECT 5.5 1.65 5.9 2.6 ;
      RECT 5.5 1.65 6.8 1.9 ;
      RECT 6.55 1.05 6.8 1.9 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 3.95 2.25 4.2 2.65 ;
      RECT 3 2.3 4.35 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 13.85 2.25 14.35 2.55 ;
      RECT 12.4 2.25 12.9 2.55 ;
      RECT 9.55 2.95 10.05 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffr_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffrn_1 0 0 ;
  SIZE 19.25 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 19.25 8.3 ;
        RECT 17.6 5.55 17.85 8.3 ;
        RECT 14.6 5.55 14.85 8.3 ;
        RECT 13.4 5.55 13.65 8.3 ;
        RECT 10.75 6.3 11 8.3 ;
        RECT 7.95 5.55 8.2 8.3 ;
        RECT 4.9 5.55 5.15 8.3 ;
        RECT 3.55 5.55 3.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 19.25 0.7 ;
        RECT 17.6 0 17.85 1.9 ;
        RECT 15.85 0 16.1 1.9 ;
        RECT 14.15 0 14.4 1.9 ;
        RECT 13.4 0 13.65 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 7.95 0 8.2 1.5 ;
        RECT 4.9 0 5.15 1.9 ;
        RECT 4 0 4.25 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 13.15 2.95 13.65 3.25 ;
      LAYER Metal2 ;
        RECT 13.15 2.9 13.65 3.3 ;
      LAYER Via1 ;
        RECT 13.27 2.97 13.53 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.4 3.6 5.9 3.9 ;
      LAYER Metal2 ;
        RECT 5.4 3.55 5.9 3.95 ;
      LAYER Via1 ;
        RECT 5.52 3.62 5.78 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 18.45 4.9 18.95 5.25 ;
        RECT 18.45 4.85 18.9 5.25 ;
        RECT 18.45 1.05 18.7 7.25 ;
      LAYER Metal2 ;
        RECT 18.45 4.9 18.95 5.2 ;
        RECT 18.5 4.85 18.9 5.25 ;
      LAYER Via1 ;
        RECT 18.57 4.92 18.83 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.75 4.25 18.2 4.55 ;
        RECT 17.85 2.15 18.1 4.55 ;
        RECT 16.75 2.15 18.1 2.4 ;
        RECT 16.75 4.25 17 7.25 ;
        RECT 16.75 1.05 17 2.4 ;
      LAYER Metal2 ;
        RECT 17.7 4.25 18.2 4.55 ;
        RECT 17.75 4.2 18.15 4.6 ;
      LAYER Via1 ;
        RECT 17.82 4.27 18.08 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  OBS
    LAYER Metal2 ;
      RECT 17 2.9 17.4 3.3 ;
      RECT 16.65 2.95 17.45 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 15.4 2.2 16 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 15.4 1 15.7 2.6 ;
      RECT 2.75 1 15.7 1.3 ;
      RECT 14.05 2.2 14.55 2.6 ;
      RECT 14.05 1.65 14.45 2.6 ;
      RECT 9.3 1.6 9.7 2 ;
      RECT 9.25 1.65 14.45 1.95 ;
      RECT 14.1 4.85 14.5 5.25 ;
      RECT 10.25 4.85 10.65 5.25 ;
      RECT 10.2 4.9 14.55 5.2 ;
      RECT 12.45 4.2 12.9 4.6 ;
      RECT 11.2 4.2 11.6 4.6 ;
      RECT 9.55 4.2 10.05 4.6 ;
      RECT 6.75 4.2 7.2 4.6 ;
      RECT 6.75 4.25 12.9 4.55 ;
      RECT 11.55 2.9 11.95 3.3 ;
      RECT 9.6 2.9 10 3.3 ;
      RECT 9.55 2.95 12.05 3.25 ;
      RECT 10.3 3.55 10.7 3.95 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 7.6 2.25 8 2.65 ;
      RECT 3.85 2.25 4.35 2.65 ;
      RECT 3.85 2.3 8.05 2.6 ;
      RECT 15.9 4.85 16.4 5.25 ;
    LAYER Via1 ;
      RECT 17.07 2.97 17.33 3.23 ;
      RECT 16.02 4.92 16.28 5.18 ;
      RECT 15.62 2.27 15.88 2.53 ;
      RECT 14.17 2.27 14.43 2.53 ;
      RECT 14.17 4.92 14.43 5.18 ;
      RECT 12.52 4.27 12.78 4.53 ;
      RECT 11.62 2.97 11.88 3.23 ;
      RECT 11.27 4.27 11.53 4.53 ;
      RECT 10.37 3.62 10.63 3.88 ;
      RECT 10.32 4.92 10.58 5.18 ;
      RECT 9.67 2.97 9.93 3.23 ;
      RECT 9.67 4.27 9.93 4.53 ;
      RECT 9.37 1.67 9.63 1.93 ;
      RECT 7.67 2.32 7.93 2.58 ;
      RECT 6.87 4.27 7.13 4.53 ;
      RECT 3.97 2.32 4.23 2.58 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 16 2.95 16.25 7.25 ;
      RECT 14.15 4.8 14.45 5.3 ;
      RECT 14.15 4.9 16.4 5.2 ;
      RECT 15 2.95 17.45 3.25 ;
      RECT 15 1.05 15.25 3.25 ;
      RECT 12.55 1.05 12.8 7.25 ;
      RECT 12.4 4.25 12.9 4.55 ;
      RECT 11.6 4.85 11.85 7.25 ;
      RECT 11.6 4.85 12.15 5.1 ;
      RECT 11.9 3.65 12.15 5.1 ;
      RECT 11.6 2.85 11.9 3.9 ;
      RECT 11.6 1.05 11.85 3.9 ;
      RECT 10.2 4.9 10.7 5.2 ;
      RECT 10.3 3.6 10.6 5.2 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 9 4.25 10.05 4.55 ;
      RECT 9 2.25 9.3 4.55 ;
      RECT 8.9 2.25 9.4 2.55 ;
      RECT 9.35 6.05 9.6 7.25 ;
      RECT 8.45 6.05 9.6 6.3 ;
      RECT 8.45 3.55 8.7 6.3 ;
      RECT 8.4 1.7 8.65 3.8 ;
      RECT 8.4 1.7 9.75 1.95 ;
      RECT 9.35 1.65 9.75 1.95 ;
      RECT 9.35 1.05 9.6 1.95 ;
      RECT 7.55 4.9 8.05 5.2 ;
      RECT 7.65 2.3 7.95 5.2 ;
      RECT 7.55 2.3 8.05 2.6 ;
      RECT 6.1 4.25 7.25 4.55 ;
      RECT 6.85 2.3 7.15 4.55 ;
      RECT 6.75 2.3 7.25 2.6 ;
      RECT 6.55 5.05 6.8 7.25 ;
      RECT 4.9 5.05 6.8 5.3 ;
      RECT 4.9 2.35 5.15 5.3 ;
      RECT 3.85 4.25 5.15 4.55 ;
      RECT 4.9 2.35 5.9 2.6 ;
      RECT 5.5 1.65 5.9 2.6 ;
      RECT 5.5 1.65 6.8 1.9 ;
      RECT 6.55 1.05 6.8 1.9 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 3.95 2.25 4.2 2.65 ;
      RECT 3 2.3 4.35 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 15.5 2.25 16 2.55 ;
      RECT 14.05 2.25 14.55 2.55 ;
      RECT 11.15 4.25 11.65 4.55 ;
      RECT 9.55 2.95 10.05 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffrn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffs_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffs_1 0 0 ;
  SIZE 15.45 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15.45 8.3 ;
        RECT 13.8 5.55 14.05 8.3 ;
        RECT 11.35 6.8 11.6 8.3 ;
        RECT 8.9 6.3 9.15 8.3 ;
        RECT 6.1 5.55 6.35 8.3 ;
        RECT 3.05 5.55 3.3 8.3 ;
        RECT 1.45 6.3 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15.45 0.7 ;
        RECT 13.8 0 14.05 1.9 ;
        RECT 10.65 0 10.9 1.9 ;
        RECT 8.9 0 9.15 1.9 ;
        RECT 6.1 0 6.35 1.5 ;
        RECT 3.05 0 3.3 1.9 ;
        RECT 2.15 0 2.4 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 9.3 4.25 9.8 4.55 ;
        RECT 7.15 4.25 8.2 4.55 ;
        RECT 7.05 2.25 7.55 2.55 ;
        RECT 7.15 2.25 7.45 4.55 ;
        RECT 4.25 4.25 5.4 4.55 ;
        RECT 4.9 2.3 5.4 2.6 ;
        RECT 5 2.3 5.3 4.55 ;
      LAYER Metal2 ;
        RECT 4.9 4.25 9.8 4.55 ;
        RECT 9.35 4.2 9.75 4.6 ;
        RECT 7.7 4.2 8.2 4.6 ;
        RECT 4.9 4.2 5.35 4.6 ;
      LAYER Via1 ;
        RECT 5.02 4.27 5.28 4.53 ;
        RECT 7.82 4.27 8.08 4.53 ;
        RECT 9.42 4.27 9.68 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 3.6 4.05 3.9 ;
      LAYER Metal2 ;
        RECT 3.55 3.55 4.05 3.95 ;
      LAYER Via1 ;
        RECT 3.67 3.62 3.93 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 14.65 4.9 15.15 5.25 ;
        RECT 14.65 4.85 15.1 5.25 ;
        RECT 14.65 1.05 14.9 7.25 ;
      LAYER Metal2 ;
        RECT 14.65 4.9 15.15 5.2 ;
        RECT 14.7 4.85 15.1 5.25 ;
      LAYER Via1 ;
        RECT 14.77 4.92 15.03 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12.95 4.25 14.4 4.55 ;
        RECT 14.05 2.15 14.3 4.55 ;
        RECT 12.95 2.15 14.3 2.4 ;
        RECT 12.95 4.25 13.2 7.25 ;
        RECT 12.95 1.05 13.2 2.4 ;
      LAYER Metal2 ;
        RECT 13.9 4.25 14.4 4.55 ;
        RECT 13.95 4.2 14.35 4.6 ;
      LAYER Via1 ;
        RECT 14.02 4.27 14.28 4.53 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.55 4.25 12.05 4.55 ;
        RECT 5.7 4.9 6.2 5.2 ;
        RECT 5.7 2.3 6.2 2.6 ;
        RECT 5.8 2.3 6.1 5.2 ;
        RECT 2.3 5.8 2.55 7.25 ;
        RECT 0.75 2.3 2.5 2.6 ;
        RECT 2.1 2.25 2.35 2.65 ;
        RECT 0.6 5.8 2.55 6.05 ;
        RECT 0.75 4.25 1.5 4.55 ;
        RECT 0.75 1.05 1 6.05 ;
        RECT 0.6 5.8 0.85 7.25 ;
      LAYER Metal2 ;
        RECT 11.55 4.2 12.05 4.6 ;
        RECT 1.1 5.55 11.95 5.85 ;
        RECT 11.65 4.2 11.95 5.85 ;
        RECT 1 4.2 1.5 4.6 ;
        RECT 1.1 4.2 1.4 5.85 ;
        RECT 2 2.3 6.2 2.6 ;
        RECT 5.75 2.25 6.15 2.65 ;
        RECT 2 2.25 2.5 2.65 ;
      LAYER Via1 ;
        RECT 1.12 4.27 1.38 4.53 ;
        RECT 2.12 2.32 2.38 2.58 ;
        RECT 5.82 2.32 6.08 2.58 ;
        RECT 11.67 4.27 11.93 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 13.2 2.9 13.6 3.3 ;
      RECT 12.85 2.95 13.65 3.25 ;
      RECT 10.55 2.2 11.05 2.6 ;
      RECT 10.55 1.65 10.95 2.6 ;
      RECT 7.45 1.6 7.85 2 ;
      RECT 7.4 1.65 10.95 1.95 ;
      RECT 10.6 4.85 11 5.25 ;
      RECT 8.4 4.85 8.8 5.25 ;
      RECT 8.35 4.9 11.05 5.2 ;
      RECT 9.7 2.9 10.1 3.3 ;
      RECT 7.75 2.9 8.15 3.3 ;
      RECT 7.7 2.95 10.2 3.25 ;
      RECT 8.45 3.55 8.85 3.95 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 12.25 4.85 12.75 5.25 ;
      RECT 2 3.55 2.5 3.95 ;
    LAYER Via1 ;
      RECT 13.27 2.97 13.53 3.23 ;
      RECT 12.37 4.92 12.63 5.18 ;
      RECT 10.67 2.27 10.93 2.53 ;
      RECT 10.67 4.92 10.93 5.18 ;
      RECT 9.77 2.97 10.03 3.23 ;
      RECT 8.52 3.62 8.78 3.88 ;
      RECT 8.47 4.92 8.73 5.18 ;
      RECT 7.82 2.97 8.08 3.23 ;
      RECT 7.52 1.67 7.78 1.93 ;
      RECT 2.12 3.62 2.38 3.88 ;
    LAYER Metal1 ;
      RECT 12.35 2.95 12.65 5.3 ;
      RECT 10.65 4.8 10.95 5.3 ;
      RECT 10.65 4.9 12.65 5.2 ;
      RECT 12.05 2.95 13.65 3.25 ;
      RECT 12.05 1.05 12.3 3.25 ;
      RECT 12.2 6.3 12.45 7.25 ;
      RECT 10.5 6.3 10.75 7.25 ;
      RECT 10.5 6.3 12.45 6.55 ;
      RECT 9.75 4.85 10 7.25 ;
      RECT 9.75 4.85 10.3 5.1 ;
      RECT 10.05 3.65 10.3 5.1 ;
      RECT 9.75 2.85 10.05 3.9 ;
      RECT 9.75 1.05 10 3.9 ;
      RECT 8.35 4.9 8.85 5.2 ;
      RECT 8.45 3.6 8.75 5.2 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 7.5 6.05 7.75 7.25 ;
      RECT 6.6 6.05 7.75 6.3 ;
      RECT 6.6 3.55 6.85 6.3 ;
      RECT 6.55 1.7 6.8 3.8 ;
      RECT 6.55 1.7 7.9 1.95 ;
      RECT 7.5 1.65 7.9 1.95 ;
      RECT 7.5 1.05 7.75 1.95 ;
      RECT 4.7 5.05 4.95 7.25 ;
      RECT 3.05 5.05 4.95 5.3 ;
      RECT 3.05 2.35 3.3 5.3 ;
      RECT 2 3.6 3.3 3.9 ;
      RECT 3.05 2.35 4.05 2.6 ;
      RECT 3.65 1.65 4.05 2.6 ;
      RECT 3.65 1.65 4.95 1.9 ;
      RECT 4.7 1.05 4.95 1.9 ;
      RECT 10.55 2.25 11.05 2.55 ;
      RECT 7.7 2.95 8.2 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffs_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsn_1 0 0 ;
  SIZE 17.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 17.2 8.3 ;
        RECT 15.5 5.55 15.75 8.3 ;
        RECT 13.05 6.8 13.3 8.3 ;
        RECT 11.45 5.55 11.7 8.3 ;
        RECT 8.9 6.3 9.15 8.3 ;
        RECT 6.1 5.55 6.35 8.3 ;
        RECT 3.05 5.55 3.3 8.3 ;
        RECT 1.45 6.3 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 17.2 0.7 ;
        RECT 15.5 0 15.75 1.9 ;
        RECT 12.35 0 12.6 1.9 ;
        RECT 11.45 0 11.7 1.9 ;
        RECT 8.9 0 9.15 1.9 ;
        RECT 6.1 0 6.35 1.5 ;
        RECT 3.05 0 3.3 1.9 ;
        RECT 2.15 0 2.4 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 11.2 2.95 11.7 3.25 ;
      LAYER Metal2 ;
        RECT 11.2 2.95 11.7 3.25 ;
        RECT 11.25 2.9 11.65 3.3 ;
      LAYER Via1 ;
        RECT 11.32 2.97 11.58 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 3.6 4.05 3.9 ;
      LAYER Metal2 ;
        RECT 3.55 3.55 4.05 3.95 ;
      LAYER Via1 ;
        RECT 3.67 3.62 3.93 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.35 4.9 16.85 5.25 ;
        RECT 16.35 4.85 16.8 5.25 ;
        RECT 16.35 1.05 16.6 7.25 ;
      LAYER Metal2 ;
        RECT 16.35 4.9 16.85 5.2 ;
        RECT 16.4 4.85 16.8 5.25 ;
      LAYER Via1 ;
        RECT 16.47 4.92 16.73 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 14.65 4.25 16.1 4.55 ;
        RECT 15.75 2.15 16 4.55 ;
        RECT 14.65 2.15 16 2.4 ;
        RECT 14.65 4.25 14.9 7.25 ;
        RECT 14.65 1.05 14.9 2.4 ;
      LAYER Metal2 ;
        RECT 15.6 4.25 16.1 4.55 ;
        RECT 15.65 4.2 16.05 4.6 ;
      LAYER Via1 ;
        RECT 15.72 4.27 15.98 4.53 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.25 4.25 13.75 4.55 ;
        RECT 5.7 4.9 6.2 5.2 ;
        RECT 5.7 2.3 6.2 2.6 ;
        RECT 5.8 2.3 6.1 5.2 ;
        RECT 2.3 5.8 2.55 7.25 ;
        RECT 0.75 2.3 2.5 2.6 ;
        RECT 2.1 2.25 2.35 2.65 ;
        RECT 0.6 5.8 2.55 6.05 ;
        RECT 0.75 4.25 1.5 4.55 ;
        RECT 0.75 1.05 1 6.05 ;
        RECT 0.6 5.8 0.85 7.25 ;
      LAYER Metal2 ;
        RECT 13.25 4.2 13.75 4.6 ;
        RECT 1.1 5.55 13.65 5.85 ;
        RECT 13.35 4.2 13.65 5.85 ;
        RECT 1 4.2 1.5 4.6 ;
        RECT 1.1 4.2 1.4 5.85 ;
        RECT 2 2.3 6.2 2.6 ;
        RECT 5.75 2.25 6.15 2.65 ;
        RECT 2 2.25 2.5 2.65 ;
      LAYER Via1 ;
        RECT 1.12 4.27 1.38 4.53 ;
        RECT 2.12 2.32 2.38 2.58 ;
        RECT 5.82 2.32 6.08 2.58 ;
        RECT 13.37 4.27 13.63 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 14.9 2.9 15.3 3.3 ;
      RECT 14.55 2.95 15.35 3.25 ;
      RECT 12.25 2.2 12.75 2.6 ;
      RECT 12.25 1.65 12.65 2.6 ;
      RECT 7.45 1.6 7.85 2 ;
      RECT 7.4 1.65 12.65 1.95 ;
      RECT 12.3 4.85 12.7 5.25 ;
      RECT 8.4 4.85 8.8 5.25 ;
      RECT 8.35 4.9 12.75 5.2 ;
      RECT 10.5 4.2 10.9 4.6 ;
      RECT 9.35 4.2 9.75 4.6 ;
      RECT 7.7 4.2 8.2 4.6 ;
      RECT 4.9 4.2 5.35 4.6 ;
      RECT 4.9 4.25 10.95 4.55 ;
      RECT 9.7 2.9 10.1 3.3 ;
      RECT 7.75 2.9 8.15 3.3 ;
      RECT 7.7 2.95 10.2 3.25 ;
      RECT 8.45 3.55 8.85 3.95 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 13.95 4.85 14.45 5.25 ;
      RECT 2 3.55 2.5 3.95 ;
    LAYER Via1 ;
      RECT 14.97 2.97 15.23 3.23 ;
      RECT 14.07 4.92 14.33 5.18 ;
      RECT 12.37 2.27 12.63 2.53 ;
      RECT 12.37 4.92 12.63 5.18 ;
      RECT 10.57 4.27 10.83 4.53 ;
      RECT 9.77 2.97 10.03 3.23 ;
      RECT 9.42 4.27 9.68 4.53 ;
      RECT 8.52 3.62 8.78 3.88 ;
      RECT 8.47 4.92 8.73 5.18 ;
      RECT 7.82 2.97 8.08 3.23 ;
      RECT 7.82 4.27 8.08 4.53 ;
      RECT 7.52 1.67 7.78 1.93 ;
      RECT 5.02 4.27 5.28 4.53 ;
      RECT 2.12 3.62 2.38 3.88 ;
    LAYER Metal1 ;
      RECT 14.05 2.95 14.35 5.3 ;
      RECT 12.35 4.8 12.65 5.3 ;
      RECT 12.35 4.9 14.35 5.2 ;
      RECT 13.75 2.95 15.35 3.25 ;
      RECT 13.75 1.05 14 3.25 ;
      RECT 13.9 6.3 14.15 7.25 ;
      RECT 12.2 6.3 12.45 7.25 ;
      RECT 12.2 6.3 14.15 6.55 ;
      RECT 10.6 1.05 10.85 7.25 ;
      RECT 10.55 1.8 10.85 5.7 ;
      RECT 10.55 4.25 10.9 4.55 ;
      RECT 9.75 4.85 10 7.25 ;
      RECT 9.75 4.85 10.3 5.1 ;
      RECT 10.05 3.65 10.3 5.1 ;
      RECT 9.75 2.85 10.05 3.9 ;
      RECT 9.75 1.05 10 3.9 ;
      RECT 8.35 4.9 8.85 5.2 ;
      RECT 8.45 3.6 8.75 5.2 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 7.15 4.25 8.2 4.55 ;
      RECT 7.15 2.25 7.45 4.55 ;
      RECT 7.05 2.25 7.55 2.55 ;
      RECT 7.5 6.05 7.75 7.25 ;
      RECT 6.6 6.05 7.75 6.3 ;
      RECT 6.6 3.55 6.85 6.3 ;
      RECT 6.55 1.7 6.8 3.8 ;
      RECT 6.55 1.7 7.9 1.95 ;
      RECT 7.5 1.65 7.9 1.95 ;
      RECT 7.5 1.05 7.75 1.95 ;
      RECT 4.25 4.25 5.4 4.55 ;
      RECT 5 2.3 5.3 4.55 ;
      RECT 4.9 2.3 5.4 2.6 ;
      RECT 4.7 5.05 4.95 7.25 ;
      RECT 3.05 5.05 4.95 5.3 ;
      RECT 3.05 2.35 3.3 5.3 ;
      RECT 2 3.6 3.3 3.9 ;
      RECT 3.05 2.35 4.05 2.6 ;
      RECT 3.65 1.65 4.05 2.6 ;
      RECT 3.65 1.65 4.95 1.9 ;
      RECT 4.7 1.05 4.95 1.9 ;
      RECT 12.25 2.25 12.75 2.55 ;
      RECT 9.3 4.25 9.8 4.55 ;
      RECT 7.7 2.95 8.2 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsr_1 0 0 ;
  SIZE 18.7 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 18.7 8.3 ;
        RECT 17.05 5.55 17.3 8.3 ;
        RECT 13.75 6.8 14 8.3 ;
        RECT 11.3 6.3 11.55 8.3 ;
        RECT 8.5 5.55 8.75 8.3 ;
        RECT 5.45 5.55 5.7 8.3 ;
        RECT 3.85 6.3 4.1 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 18.7 0.7 ;
        RECT 17.05 0 17.3 1.9 ;
        RECT 15.3 0 15.55 1.9 ;
        RECT 13.05 0 13.3 1.9 ;
        RECT 11.3 0 11.55 1.9 ;
        RECT 8.5 0 8.75 1.5 ;
        RECT 5.45 0 5.7 1.9 ;
        RECT 4.55 0 4.8 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 11.7 4.25 12.2 4.55 ;
        RECT 9.55 4.25 10.6 4.55 ;
        RECT 9.45 2.25 9.95 2.55 ;
        RECT 9.55 2.25 9.85 4.55 ;
        RECT 6.65 4.25 7.8 4.55 ;
        RECT 7.3 2.3 7.8 2.6 ;
        RECT 7.4 2.3 7.7 4.55 ;
      LAYER Metal2 ;
        RECT 7.3 4.25 12.2 4.55 ;
        RECT 11.75 4.2 12.15 4.6 ;
        RECT 10.1 4.2 10.6 4.6 ;
        RECT 7.3 4.2 7.75 4.6 ;
      LAYER Via1 ;
        RECT 7.42 4.27 7.68 4.53 ;
        RECT 10.22 4.27 10.48 4.53 ;
        RECT 11.82 4.27 12.08 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 3.6 6.45 3.9 ;
      LAYER Metal2 ;
        RECT 5.95 3.55 6.45 3.95 ;
      LAYER Via1 ;
        RECT 6.07 3.62 6.33 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17.9 4.9 18.4 5.25 ;
        RECT 17.9 4.85 18.35 5.25 ;
        RECT 17.9 1.05 18.15 7.25 ;
      LAYER Metal2 ;
        RECT 17.9 4.9 18.4 5.2 ;
        RECT 17.95 4.85 18.35 5.25 ;
      LAYER Via1 ;
        RECT 18.02 4.92 18.28 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.2 4.25 17.65 4.55 ;
        RECT 17.3 2.15 17.55 4.55 ;
        RECT 16.2 2.15 17.55 2.4 ;
        RECT 16.2 4.25 16.45 7.25 ;
        RECT 16.2 1.05 16.45 2.4 ;
      LAYER Metal2 ;
        RECT 17.15 4.25 17.65 4.55 ;
        RECT 17.2 4.2 17.6 4.6 ;
      LAYER Via1 ;
        RECT 17.27 4.27 17.53 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.95 4.25 14.45 4.55 ;
        RECT 3.4 4.25 3.9 4.55 ;
      LAYER Metal2 ;
        RECT 13.95 4.2 14.45 4.6 ;
        RECT 3.5 5.55 14.35 5.85 ;
        RECT 14.05 4.2 14.35 5.85 ;
        RECT 3.4 4.2 3.9 4.6 ;
        RECT 3.5 4.2 3.8 5.85 ;
      LAYER Via1 ;
        RECT 3.52 4.27 3.78 4.53 ;
        RECT 14.07 4.27 14.33 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 16.45 2.9 16.85 3.3 ;
      RECT 16.1 2.95 16.9 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 14.85 2.2 15.45 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 14.85 1 15.15 2.6 ;
      RECT 2.75 1 15.15 1.3 ;
      RECT 12.95 2.2 13.45 2.6 ;
      RECT 12.95 1.65 13.35 2.6 ;
      RECT 9.85 1.6 10.25 2 ;
      RECT 9.8 1.65 13.35 1.95 ;
      RECT 13 4.85 13.4 5.25 ;
      RECT 10.8 4.85 11.2 5.25 ;
      RECT 10.75 4.9 13.45 5.2 ;
      RECT 12.1 2.9 12.5 3.3 ;
      RECT 10.15 2.9 10.55 3.3 ;
      RECT 10.1 2.95 12.6 3.25 ;
      RECT 10.85 3.55 11.25 3.95 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 8.15 2.25 8.55 2.65 ;
      RECT 4.4 2.25 4.9 2.65 ;
      RECT 4.4 2.3 8.6 2.6 ;
      RECT 15.35 4.85 15.85 5.25 ;
      RECT 4.4 3.55 4.9 3.95 ;
    LAYER Via1 ;
      RECT 16.52 2.97 16.78 3.23 ;
      RECT 15.47 4.92 15.73 5.18 ;
      RECT 15.07 2.27 15.33 2.53 ;
      RECT 13.07 2.27 13.33 2.53 ;
      RECT 13.07 4.92 13.33 5.18 ;
      RECT 12.17 2.97 12.43 3.23 ;
      RECT 10.92 3.62 11.18 3.88 ;
      RECT 10.87 4.92 11.13 5.18 ;
      RECT 10.22 2.97 10.48 3.23 ;
      RECT 9.92 1.67 10.18 1.93 ;
      RECT 8.22 2.32 8.48 2.58 ;
      RECT 4.52 2.32 4.78 2.58 ;
      RECT 4.52 3.62 4.78 3.88 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 15.45 2.95 15.7 7.25 ;
      RECT 13.05 4.8 13.35 5.3 ;
      RECT 13.05 4.9 15.85 5.2 ;
      RECT 14.45 2.95 16.9 3.25 ;
      RECT 14.45 1.05 14.7 3.25 ;
      RECT 14.6 6.3 14.85 7.25 ;
      RECT 12.9 6.3 13.15 7.25 ;
      RECT 12.9 6.3 14.85 6.55 ;
      RECT 12.15 4.85 12.4 7.25 ;
      RECT 12.15 4.85 12.7 5.1 ;
      RECT 12.45 3.65 12.7 5.1 ;
      RECT 12.15 2.85 12.45 3.9 ;
      RECT 12.15 1.05 12.4 3.9 ;
      RECT 10.75 4.9 11.25 5.2 ;
      RECT 10.85 3.6 11.15 5.2 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 9.9 6.05 10.15 7.25 ;
      RECT 9 6.05 10.15 6.3 ;
      RECT 9 3.55 9.25 6.3 ;
      RECT 8.95 1.7 9.2 3.8 ;
      RECT 8.95 1.7 10.3 1.95 ;
      RECT 9.9 1.65 10.3 1.95 ;
      RECT 9.9 1.05 10.15 1.95 ;
      RECT 8.1 4.9 8.6 5.2 ;
      RECT 8.2 2.3 8.5 5.2 ;
      RECT 8.1 2.3 8.6 2.6 ;
      RECT 7.1 5.05 7.35 7.25 ;
      RECT 5.45 5.05 7.35 5.3 ;
      RECT 5.45 2.35 5.7 5.3 ;
      RECT 4.4 3.6 5.7 3.9 ;
      RECT 5.45 2.35 6.45 2.6 ;
      RECT 6.05 1.65 6.45 2.6 ;
      RECT 6.05 1.65 7.35 1.9 ;
      RECT 7.1 1.05 7.35 1.9 ;
      RECT 4.7 5.8 4.95 7.25 ;
      RECT 3 5.8 3.25 7.25 ;
      RECT 3 5.8 4.95 6.05 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 4.5 2.25 4.75 2.65 ;
      RECT 3.15 2.3 4.9 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 14.95 2.25 15.45 2.55 ;
      RECT 12.95 2.25 13.45 2.55 ;
      RECT 10.1 2.95 10.6 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsr_1

MACRO gf180mcu_osu_sc_gp12t3v3__dffsrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsrn_1 0 0 ;
  SIZE 20.45 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 20.45 8.3 ;
        RECT 18.8 5.55 19.05 8.3 ;
        RECT 15.5 6.8 15.75 8.3 ;
        RECT 13.9 5.55 14.15 8.3 ;
        RECT 11.3 6.3 11.55 8.3 ;
        RECT 8.5 5.55 8.75 8.3 ;
        RECT 5.45 5.55 5.7 8.3 ;
        RECT 3.85 6.3 4.1 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 20.45 0.7 ;
        RECT 18.8 0 19.05 1.9 ;
        RECT 17.05 0 17.3 1.9 ;
        RECT 14.8 0 15.05 1.9 ;
        RECT 13.9 0 14.15 1.9 ;
        RECT 11.3 0 11.55 1.9 ;
        RECT 8.5 0 8.75 1.5 ;
        RECT 5.45 0 5.7 1.9 ;
        RECT 4.55 0 4.8 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 13.65 2.95 14.15 3.25 ;
      LAYER Metal2 ;
        RECT 13.65 2.9 14.15 3.3 ;
      LAYER Via1 ;
        RECT 13.77 2.97 14.03 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 3.6 6.45 3.9 ;
      LAYER Metal2 ;
        RECT 5.95 3.55 6.45 3.95 ;
      LAYER Via1 ;
        RECT 6.07 3.62 6.33 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 19.65 4.9 20.15 5.25 ;
        RECT 19.65 4.85 20.1 5.25 ;
        RECT 19.65 1.05 19.9 7.25 ;
      LAYER Metal2 ;
        RECT 19.65 4.9 20.15 5.2 ;
        RECT 19.7 4.85 20.1 5.25 ;
      LAYER Via1 ;
        RECT 19.77 4.92 20.03 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17.95 4.25 19.4 4.55 ;
        RECT 19.05 2.15 19.3 4.55 ;
        RECT 17.95 2.15 19.3 2.4 ;
        RECT 17.95 4.25 18.2 7.25 ;
        RECT 17.95 1.05 18.2 2.4 ;
      LAYER Metal2 ;
        RECT 18.9 4.25 19.4 4.55 ;
        RECT 18.95 4.2 19.35 4.6 ;
      LAYER Via1 ;
        RECT 19.02 4.27 19.28 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15.7 4.25 16.2 4.55 ;
        RECT 3.4 4.25 3.9 4.55 ;
      LAYER Metal2 ;
        RECT 15.7 4.2 16.2 4.6 ;
        RECT 3.5 5.55 16.1 5.85 ;
        RECT 15.8 4.2 16.1 5.85 ;
        RECT 3.4 4.2 3.9 4.6 ;
        RECT 3.5 4.2 3.8 5.85 ;
      LAYER Via1 ;
        RECT 3.52 4.27 3.78 4.53 ;
        RECT 15.82 4.27 16.08 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 18.2 2.9 18.6 3.3 ;
      RECT 17.85 2.95 18.65 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 16.6 2.2 17.2 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 16.6 1 16.9 2.6 ;
      RECT 2.75 1 16.9 1.3 ;
      RECT 14.7 2.2 15.2 2.6 ;
      RECT 14.7 1.65 15.1 2.6 ;
      RECT 9.85 1.6 10.25 2 ;
      RECT 9.8 1.65 15.1 1.95 ;
      RECT 14.75 4.85 15.15 5.25 ;
      RECT 10.8 4.85 11.2 5.25 ;
      RECT 10.75 4.9 15.2 5.2 ;
      RECT 12.95 4.2 13.4 4.6 ;
      RECT 11.75 4.2 12.15 4.6 ;
      RECT 10.1 4.2 10.6 4.6 ;
      RECT 7.3 4.2 7.75 4.6 ;
      RECT 7.3 4.25 13.4 4.55 ;
      RECT 12.1 2.9 12.5 3.3 ;
      RECT 10.15 2.9 10.55 3.3 ;
      RECT 10.1 2.95 12.6 3.25 ;
      RECT 10.85 3.55 11.25 3.95 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 8.15 2.25 8.55 2.65 ;
      RECT 4.4 2.25 4.9 2.65 ;
      RECT 4.4 2.3 8.6 2.6 ;
      RECT 17.1 4.85 17.6 5.25 ;
      RECT 4.4 3.55 4.9 3.95 ;
    LAYER Via1 ;
      RECT 18.27 2.97 18.53 3.23 ;
      RECT 17.22 4.92 17.48 5.18 ;
      RECT 16.82 2.27 17.08 2.53 ;
      RECT 14.82 2.27 15.08 2.53 ;
      RECT 14.82 4.92 15.08 5.18 ;
      RECT 13.02 4.27 13.28 4.53 ;
      RECT 12.17 2.97 12.43 3.23 ;
      RECT 11.82 4.27 12.08 4.53 ;
      RECT 10.92 3.62 11.18 3.88 ;
      RECT 10.87 4.92 11.13 5.18 ;
      RECT 10.22 2.97 10.48 3.23 ;
      RECT 10.22 4.27 10.48 4.53 ;
      RECT 9.92 1.67 10.18 1.93 ;
      RECT 8.22 2.32 8.48 2.58 ;
      RECT 7.42 4.27 7.68 4.53 ;
      RECT 4.52 2.32 4.78 2.58 ;
      RECT 4.52 3.62 4.78 3.88 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 17.2 2.95 17.45 7.25 ;
      RECT 14.8 4.8 15.1 5.3 ;
      RECT 14.8 4.9 17.6 5.2 ;
      RECT 16.2 2.95 18.65 3.25 ;
      RECT 16.2 1.05 16.45 3.25 ;
      RECT 16.35 6.3 16.6 7.25 ;
      RECT 14.65 6.3 14.9 7.25 ;
      RECT 14.65 6.3 16.6 6.55 ;
      RECT 13.05 1.05 13.3 7.25 ;
      RECT 13 1.8 13.3 5.65 ;
      RECT 12.95 4.25 13.4 4.55 ;
      RECT 12.15 4.85 12.4 7.25 ;
      RECT 12.15 4.85 12.7 5.1 ;
      RECT 12.45 3.65 12.7 5.1 ;
      RECT 12.15 2.85 12.45 3.9 ;
      RECT 12.15 1.05 12.4 3.9 ;
      RECT 10.75 4.9 11.25 5.2 ;
      RECT 10.85 3.6 11.15 5.2 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 9.55 4.25 10.6 4.55 ;
      RECT 9.55 2.25 9.85 4.55 ;
      RECT 9.45 2.25 9.95 2.55 ;
      RECT 9.9 6.05 10.15 7.25 ;
      RECT 9 6.05 10.15 6.3 ;
      RECT 9 3.55 9.25 6.3 ;
      RECT 8.95 1.7 9.2 3.8 ;
      RECT 8.95 1.7 10.3 1.95 ;
      RECT 9.9 1.65 10.3 1.95 ;
      RECT 9.9 1.05 10.15 1.95 ;
      RECT 8.1 4.9 8.6 5.2 ;
      RECT 8.2 2.3 8.5 5.2 ;
      RECT 8.1 2.3 8.6 2.6 ;
      RECT 6.65 4.25 7.8 4.55 ;
      RECT 7.4 2.3 7.7 4.55 ;
      RECT 7.3 2.3 7.8 2.6 ;
      RECT 7.1 5.05 7.35 7.25 ;
      RECT 5.45 5.05 7.35 5.3 ;
      RECT 5.45 2.35 5.7 5.3 ;
      RECT 4.4 3.6 5.7 3.9 ;
      RECT 5.45 2.35 6.45 2.6 ;
      RECT 6.05 1.65 6.45 2.6 ;
      RECT 6.05 1.65 7.35 1.9 ;
      RECT 7.1 1.05 7.35 1.9 ;
      RECT 4.7 5.8 4.95 7.25 ;
      RECT 3 5.8 3.25 7.25 ;
      RECT 3 5.8 4.95 6.05 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 4.5 2.25 4.75 2.65 ;
      RECT 3.15 2.3 4.9 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 16.7 2.25 17.2 2.55 ;
      RECT 14.7 2.25 15.2 2.55 ;
      RECT 11.7 4.25 12.2 4.55 ;
      RECT 10.1 2.95 10.6 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsrn_1

MACRO gf180mcu_osu_sc_gp12t3v3__dlat_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlat_1 0 0 ;
  SIZE 9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal2 ;
        RECT 5.2 4.2 5.7 4.6 ;
        RECT 3.45 4.25 5.7 4.55 ;
        RECT 3.5 4.2 3.9 4.6 ;
      LAYER Metal1 ;
        RECT 5.2 4.25 5.7 4.55 ;
        RECT 3.45 4.25 3.95 4.55 ;
      LAYER Via1 ;
        RECT 3.57 4.27 3.83 4.53 ;
        RECT 5.32 4.27 5.58 4.53 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 9 8.3 ;
        RECT 7.3 5.55 7.55 8.3 ;
        RECT 4.85 5.55 5.1 8.3 ;
        RECT 1.45 6.35 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 9 0.7 ;
        RECT 7.3 0 7.55 1.9 ;
        RECT 4.7 0 5.1 1.9 ;
        RECT 1.45 0 1.85 1.9 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.85 4.2 2.35 4.6 ;
      LAYER Metal1 ;
        RECT 1.85 4.25 2.35 4.55 ;
      LAYER Via1 ;
        RECT 1.97 4.27 2.23 4.53 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.15 4.9 8.65 5.2 ;
        RECT 8.2 4.85 8.6 5.25 ;
      LAYER Metal1 ;
        RECT 8.15 4.9 8.65 5.2 ;
        RECT 8.15 4.85 8.55 5.25 ;
        RECT 8.15 1.05 8.4 7.25 ;
      LAYER Via1 ;
        RECT 8.27 4.92 8.53 5.18 ;
    END
  END Q
  OBS
    LAYER Metal2 ;
      RECT 6.75 3.55 7.25 3.95 ;
      RECT 4.55 3.55 4.95 3.95 ;
      RECT 0.35 3.55 0.85 3.95 ;
      RECT 0.35 3.6 7.25 3.9 ;
      RECT 6.5 4.85 6.9 5.25 ;
      RECT 6.45 4.9 6.95 5.2 ;
    LAYER Via1 ;
      RECT 6.87 3.62 7.13 3.88 ;
      RECT 6.57 4.92 6.83 5.18 ;
      RECT 4.62 3.62 4.88 3.88 ;
      RECT 0.47 3.62 0.73 3.88 ;
    LAYER Metal1 ;
      RECT 6.45 4.85 6.7 7.25 ;
      RECT 6.45 4.85 6.85 5.4 ;
      RECT 6.45 4.9 6.95 5.2 ;
      RECT 6.45 4.9 7.8 5.15 ;
      RECT 7.5 2.15 7.8 5.15 ;
      RECT 6.45 2.15 7.8 2.4 ;
      RECT 6.45 1.05 6.7 2.4 ;
      RECT 5.7 5.35 5.95 7.25 ;
      RECT 5.95 2.05 6.2 5.6 ;
      RECT 2.6 4.8 3.1 5.1 ;
      RECT 2.7 2.65 3 5.1 ;
      RECT 2.7 2.65 6.2 2.95 ;
      RECT 5.7 1.05 5.95 2.3 ;
      RECT 3.15 5.55 3.4 7.25 ;
      RECT 1.15 5.55 3.4 5.8 ;
      RECT 1.15 2.15 1.4 5.8 ;
      RECT 1.1 4.25 1.55 4.55 ;
      RECT 1.15 2.15 3.4 2.4 ;
      RECT 3.15 1.05 3.4 2.4 ;
      RECT 0.6 1.05 0.85 7.25 ;
      RECT 0.5 3.55 0.85 3.95 ;
      RECT 0.35 3.6 0.85 3.9 ;
      RECT 0.45 3.55 0.85 3.9 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 4.5 3.6 5 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlat_1

MACRO gf180mcu_osu_sc_gp12t3v3__dlatn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlatn_1 0 0 ;
  SIZE 10.7 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 10.7 8.3 ;
        RECT 9 5.55 9.25 8.3 ;
        RECT 7.4 5.55 7.65 8.3 ;
        RECT 4.85 5.55 5.1 8.3 ;
        RECT 1.45 6.35 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 10.7 0.7 ;
        RECT 9 0 9.25 1.9 ;
        RECT 7.4 0 7.65 1.9 ;
        RECT 4.7 0 5.1 1.9 ;
        RECT 1.45 0 1.85 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 7.05 2.65 7.55 2.95 ;
      LAYER Metal2 ;
        RECT 7.05 2.6 7.55 3 ;
      LAYER Via1 ;
        RECT 7.17 2.67 7.43 2.93 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.85 4.25 2.35 4.55 ;
      LAYER Metal2 ;
        RECT 1.85 4.2 2.35 4.6 ;
      LAYER Via1 ;
        RECT 1.97 4.27 2.23 4.53 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.85 4.9 10.35 5.2 ;
        RECT 9.85 4.85 10.25 5.25 ;
        RECT 9.85 1.05 10.1 7.25 ;
      LAYER Metal2 ;
        RECT 9.85 4.9 10.35 5.2 ;
        RECT 9.9 4.85 10.3 5.25 ;
      LAYER Via1 ;
        RECT 9.97 4.92 10.23 5.18 ;
    END
  END Q
  OBS
    LAYER Metal2 ;
      RECT 8.45 3.55 8.95 3.95 ;
      RECT 4.55 3.55 4.95 3.95 ;
      RECT 0.35 3.55 0.85 3.95 ;
      RECT 0.35 3.6 8.95 3.9 ;
      RECT 8.2 4.85 8.6 5.25 ;
      RECT 8.15 4.9 8.65 5.2 ;
      RECT 6.45 4.2 6.95 4.6 ;
      RECT 5.2 4.2 5.7 4.6 ;
      RECT 3.5 4.2 3.9 4.6 ;
      RECT 3.45 4.25 6.95 4.55 ;
    LAYER Via1 ;
      RECT 8.57 3.62 8.83 3.88 ;
      RECT 8.27 4.92 8.53 5.18 ;
      RECT 6.57 4.27 6.83 4.53 ;
      RECT 5.32 4.27 5.58 4.53 ;
      RECT 4.62 3.62 4.88 3.88 ;
      RECT 3.57 4.27 3.83 4.53 ;
      RECT 0.47 3.62 0.73 3.88 ;
    LAYER Metal1 ;
      RECT 8.15 4.85 8.4 7.25 ;
      RECT 8.15 4.85 8.55 5.4 ;
      RECT 8.15 4.9 8.65 5.2 ;
      RECT 8.15 4.9 9.5 5.15 ;
      RECT 9.2 2.15 9.5 5.15 ;
      RECT 8.15 2.15 9.5 2.4 ;
      RECT 8.15 1.05 8.4 2.4 ;
      RECT 6.55 1.05 6.8 7.25 ;
      RECT 6.55 4.2 6.95 4.6 ;
      RECT 6.45 4.25 6.95 4.55 ;
      RECT 5.7 5.35 5.95 7.25 ;
      RECT 5.95 2.05 6.2 5.6 ;
      RECT 2.6 4.8 3.1 5.1 ;
      RECT 2.7 2.65 3 5.1 ;
      RECT 2.7 2.65 6.2 2.95 ;
      RECT 5.7 1.05 5.95 2.3 ;
      RECT 3.15 5.55 3.4 7.25 ;
      RECT 1.15 5.55 3.4 5.8 ;
      RECT 1.15 2.15 1.4 5.8 ;
      RECT 1.1 4.25 1.55 4.55 ;
      RECT 1.15 2.15 3.4 2.4 ;
      RECT 3.15 1.05 3.4 2.4 ;
      RECT 0.6 1.05 0.85 7.25 ;
      RECT 0.5 3.55 0.85 3.95 ;
      RECT 0.35 3.6 0.85 3.9 ;
      RECT 0.45 3.55 0.85 3.9 ;
      RECT 8.45 3.6 8.95 3.9 ;
      RECT 5.2 4.25 5.7 4.55 ;
      RECT 4.5 3.6 5 3.9 ;
      RECT 3.45 4.25 3.95 4.55 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlatn_1

MACRO gf180mcu_osu_sc_gp12t3v3__fill_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_1 0 0 ;
  SIZE 0.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 0.1 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 0.1 0.7 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_1

MACRO gf180mcu_osu_sc_gp12t3v3__fill_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_16 0 0 ;
  SIZE 1.6 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 1.6 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 1.6 0.7 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_16

MACRO gf180mcu_osu_sc_gp12t3v3__fill_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_2 0 0 ;
  SIZE 0.2 BY 8.2 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 0.2 8.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 0.2 0.7 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_2

MACRO gf180mcu_osu_sc_gp12t3v3__fill_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_4 0 0 ;
  SIZE 0.4 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 0.4 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 0.4 0.7 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_4

MACRO gf180mcu_osu_sc_gp12t3v3__fill_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__fill_8 0 0 ;
  SIZE 0.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 0.8 0.7 ;
    END
  END VSS
END gf180mcu_osu_sc_gp12t3v3__fill_8

MACRO gf180mcu_osu_sc_gp12t3v3__inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_1 0 0 ;
  SIZE 2.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.2 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.2 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 3.6 1.8 3.9 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 1.3 3.55 1.8 3.95 ;
      LAYER Via1 ;
        RECT 1.42 3.62 1.68 3.88 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_1

MACRO gf180mcu_osu_sc_gp12t3v3__inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_16 0 0 ;
  SIZE 15 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15 8.3 ;
        RECT 14.15 5.55 14.4 8.3 ;
        RECT 12.45 5.55 12.7 8.3 ;
        RECT 10.75 5.55 11 8.3 ;
        RECT 9.05 5.55 9.3 8.3 ;
        RECT 7.35 5.55 7.6 8.3 ;
        RECT 5.65 5.55 5.9 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15 0.7 ;
        RECT 14.15 0 14.4 1.9 ;
        RECT 12.45 0 12.7 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 9.05 0 9.3 1.9 ;
        RECT 7.35 0 7.6 1.9 ;
        RECT 5.65 0 5.9 1.9 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.3 1.05 13.55 7.25 ;
        RECT 1.4 4.55 13.55 4.8 ;
        RECT 13.15 4.2 13.55 4.8 ;
        RECT 1.4 2.15 13.55 2.4 ;
        RECT 11.6 1.05 11.85 7.25 ;
        RECT 9.9 1.05 10.15 7.25 ;
        RECT 8.2 1.05 8.45 7.25 ;
        RECT 6.5 1.05 6.75 7.25 ;
        RECT 4.8 1.05 5.05 7.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 13.15 4.2 13.65 4.6 ;
      LAYER Via1 ;
        RECT 13.27 4.27 13.53 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_16

MACRO gf180mcu_osu_sc_gp12t3v3__inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_2 0 0 ;
  SIZE 3.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.2 8.3 ;
        RECT 2.3 5.55 2.55 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.2 0.7 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 3.6 1.15 3.9 ;
      LAYER Metal2 ;
        RECT 0.65 3.55 1.15 3.95 ;
      LAYER Via1 ;
        RECT 0.77 3.62 1.03 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.4 4.25 2 4.55 ;
        RECT 1.4 4.1 1.85 4.65 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 1.5 4.2 2 4.6 ;
      LAYER Via1 ;
        RECT 1.62 4.27 1.88 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_2

MACRO gf180mcu_osu_sc_gp12t3v3__inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_4 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 4.55 3.35 4.8 ;
        RECT 2.95 4.2 3.35 4.8 ;
        RECT 1.4 2.15 3.35 2.4 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 2.95 4.2 3.45 4.6 ;
      LAYER Via1 ;
        RECT 3.07 4.27 3.33 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_4

MACRO gf180mcu_osu_sc_gp12t3v3__inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__inv_8 0 0 ;
  SIZE 8.15 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 8.15 8.3 ;
        RECT 7.35 5.55 7.6 8.3 ;
        RECT 5.65 5.55 5.9 8.3 ;
        RECT 3.95 5.55 4.2 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 8.15 0.7 ;
        RECT 7.35 0 7.6 1.9 ;
        RECT 5.65 0 5.9 1.9 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 3.6 0.9 3.9 ;
      LAYER Metal2 ;
        RECT 0.4 3.55 0.9 3.95 ;
      LAYER Via1 ;
        RECT 0.52 3.62 0.78 3.88 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.5 1.05 6.75 7.25 ;
        RECT 1.4 4.55 6.75 4.8 ;
        RECT 6.35 4.2 6.75 4.8 ;
        RECT 1.4 2.15 6.75 2.4 ;
        RECT 4.8 1.05 5.05 7.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
        RECT 1.4 1.05 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 6.35 4.2 6.85 4.6 ;
      LAYER Via1 ;
        RECT 6.47 4.27 6.73 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__inv_8

MACRO gf180mcu_osu_sc_gp12t3v3__lshifdown
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifdown 0 0 ;
  SIZE 5.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 7.6 5.2 8.3 ;
        RECT 3.45 5.55 3.75 8.3 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.3 8.3 ;
        RECT 0.55 5.55 0.85 8.3 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.2 0.7 ;
        RECT 3.45 0 3.75 1.9 ;
        RECT 0.55 0 0.85 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.3 4.25 4.7 4.55 ;
        RECT 4.35 1.05 4.65 7.25 ;
      LAYER Metal2 ;
        RECT 4.25 4.2 4.75 4.6 ;
      LAYER Via1 ;
        RECT 4.37 4.27 4.63 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 3.5 4.85 4 5.25 ;
      RECT 1.35 4.85 1.85 5.25 ;
      RECT 1.35 4.9 4 5.2 ;
    LAYER Via1 ;
      RECT 3.62 4.92 3.88 5.18 ;
      RECT 1.47 4.92 1.73 5.18 ;
    LAYER Metal1 ;
      RECT 1.45 1.05 1.75 7.25 ;
      RECT 1.35 4.9 1.85 5.2 ;
      RECT 3.5 4.9 4 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifdown

MACRO gf180mcu_osu_sc_gp12t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifup 0 0 ;
  SIZE 7.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.3 8.3 ;
        RECT 0.55 5.55 0.85 8.3 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 7.6 7.8 8.3 ;
        RECT 6.05 5.55 6.35 8.3 ;
        RECT 4.35 5.55 4.65 8.3 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 7.8 0.7 ;
        RECT 6.05 0 6.35 1.9 ;
        RECT 4.35 0 4.65 1.9 ;
        RECT 0.55 0 0.85 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4 2.3 4.5 2.6 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 4 2.25 4.5 2.65 ;
        RECT 0.6 2.3 4.5 2.6 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
        RECT 4.12 2.32 4.38 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.9 4.25 7.3 4.55 ;
        RECT 6.95 1.05 7.25 7.25 ;
      LAYER Metal2 ;
        RECT 6.85 4.2 7.35 4.6 ;
      LAYER Via1 ;
        RECT 6.97 4.27 7.23 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 6.1 4.85 6.6 5.25 ;
      RECT 4.55 4.85 4.95 5.25 ;
      RECT 4.5 4.9 6.6 5.2 ;
      RECT 4.5 2.95 5 3.35 ;
      RECT 1.35 2.95 1.85 3.35 ;
      RECT 1.35 3 5 3.3 ;
    LAYER Via1 ;
      RECT 6.22 4.92 6.48 5.18 ;
      RECT 4.62 3.02 4.88 3.28 ;
      RECT 4.62 4.92 4.88 5.18 ;
      RECT 1.47 3.02 1.73 3.28 ;
    LAYER Metal1 ;
      RECT 5.25 1.05 5.55 7.25 ;
      RECT 4.8 4.1 5.55 4.55 ;
      RECT 3.45 1.05 3.75 7.25 ;
      RECT 4.55 4.85 5 5.3 ;
      RECT 3.45 4.9 5 5.2 ;
      RECT 1.45 1.05 1.75 7.25 ;
      RECT 1.35 3 1.85 3.3 ;
      RECT 6.1 4.9 6.6 5.2 ;
      RECT 4.5 3 5 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifup

MACRO gf180mcu_osu_sc_gp12t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__mux2_1 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 3.55 2.85 3.95 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.35 3.55 2.85 3.95 ;
      LAYER Via1 ;
        RECT 2.47 3.62 2.73 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.75 4.2 4.25 4.6 ;
        RECT 3.95 1.05 4.2 7.25 ;
      LAYER Metal2 ;
        RECT 3.75 4.2 4.25 4.6 ;
      LAYER Via1 ;
        RECT 3.87 4.27 4.13 4.53 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 2.95 1.05 3.25 ;
      LAYER Metal2 ;
        RECT 0.55 2.9 1.05 3.3 ;
      LAYER Via1 ;
        RECT 0.67 2.97 0.93 3.23 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 4.85 3.5 5.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
      LAYER Metal2 ;
        RECT 3 4.85 3.5 5.25 ;
      LAYER Via1 ;
        RECT 3.12 4.92 3.38 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.4 4.25 2 4.55 ;
      RECT 1.4 2.3 2 2.6 ;
  END
END gf180mcu_osu_sc_gp12t3v3__mux2_1

MACRO gf180mcu_osu_sc_gp12t3v3__nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nand2_1 0 0 ;
  SIZE 3.1 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.1 8.3 ;
        RECT 2.25 5.55 2.5 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.1 0.7 ;
        RECT 2.1 0 2.35 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.55 1.1 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.9 2.95 2.4 3.25 ;
      LAYER Metal2 ;
        RECT 1.9 2.9 2.4 3.3 ;
      LAYER Via1 ;
        RECT 2.02 2.97 2.28 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 4.25 1.8 4.55 ;
        RECT 1.4 2 1.65 7.25 ;
        RECT 0.7 2 1.65 2.25 ;
        RECT 0.7 1.05 0.95 2.25 ;
      LAYER Metal2 ;
        RECT 1.3 4.2 1.8 4.6 ;
      LAYER Via1 ;
        RECT 1.42 4.27 1.68 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__nand2_1

MACRO gf180mcu_osu_sc_gp12t3v3__nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor2_1 0 0 ;
  SIZE 2.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.8 0.7 ;
        RECT 2.1 0 2.35 1.9 ;
        RECT 0.4 0 0.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 3.6 0.95 3.9 ;
      LAYER Metal2 ;
        RECT 0.45 3.55 0.95 3.95 ;
      LAYER Via1 ;
        RECT 0.57 3.62 0.83 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.85 2.95 2.35 3.25 ;
      LAYER Metal2 ;
        RECT 1.85 2.9 2.35 3.3 ;
      LAYER Via1 ;
        RECT 1.97 2.97 2.23 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 4.85 2.2 7.25 ;
        RECT 1.25 4.85 2.2 5.1 ;
        RECT 1.15 4.25 1.65 4.55 ;
        RECT 1.25 1.05 1.5 5.1 ;
      LAYER Metal2 ;
        RECT 1.15 4.2 1.65 4.6 ;
      LAYER Via1 ;
        RECT 1.27 4.27 1.53 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__nor2_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai21_1 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 2.95 5.55 3.2 8.3 ;
        RECT 0.65 5.55 0.9 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 1.35 0 1.6 1.6 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 3.6 0.95 3.9 ;
      LAYER Metal2 ;
        RECT 0.45 3.55 0.95 3.95 ;
      LAYER Via1 ;
        RECT 0.57 3.62 0.83 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 4.25 1.95 4.55 ;
      LAYER Metal2 ;
        RECT 1.45 4.2 1.95 4.6 ;
      LAYER Via1 ;
        RECT 1.57 4.27 1.83 4.53 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 3.6 2.7 3.9 ;
      LAYER Metal2 ;
        RECT 2.2 3.55 2.7 3.95 ;
      LAYER Via1 ;
        RECT 2.32 3.62 2.58 3.88 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 4.9 3.35 5.2 ;
        RECT 3.05 1.05 3.3 2.6 ;
        RECT 2.95 2.35 3.2 5.2 ;
        RECT 2.1 4.9 2.35 7.25 ;
      LAYER Metal2 ;
        RECT 2.85 4.85 3.35 5.25 ;
      LAYER Via1 ;
        RECT 2.97 4.92 3.23 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.5 1.85 2.45 2.1 ;
      RECT 2.2 1.05 2.45 2.1 ;
      RECT 0.5 1.05 0.75 2.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai21_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai22_1 0 0 ;
  SIZE 5.3 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.3 8.3 ;
        RECT 3.5 5.55 3.75 8.3 ;
        RECT 0.65 5.55 0.9 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.3 0.7 ;
        RECT 1.35 0 1.6 1.7 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 3.6 0.95 3.9 ;
      LAYER Metal2 ;
        RECT 0.45 3.55 0.95 3.95 ;
      LAYER Via1 ;
        RECT 0.57 3.62 0.83 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 4.25 1.95 4.55 ;
      LAYER Metal2 ;
        RECT 1.45 4.2 1.95 4.6 ;
      LAYER Via1 ;
        RECT 1.57 4.27 1.83 4.53 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 3.6 2.7 3.9 ;
      LAYER Metal2 ;
        RECT 2.2 3.55 2.7 3.95 ;
      LAYER Via1 ;
        RECT 2.32 3.62 2.58 3.88 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.15 3.6 3.65 3.9 ;
      LAYER Metal2 ;
        RECT 3.15 3.55 3.65 3.95 ;
      LAYER Via1 ;
        RECT 3.27 3.62 3.53 3.88 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.3 4.25 4.8 4.55 ;
        RECT 4.4 0.95 4.7 1.45 ;
        RECT 2.1 5 4.65 5.3 ;
        RECT 4.4 0.95 4.65 5.3 ;
        RECT 2.1 5 2.35 7.25 ;
        RECT 2.95 1 3.45 1.3 ;
        RECT 3.05 1 3.3 1.7 ;
      LAYER Metal2 ;
        RECT 4.3 4.2 4.8 4.6 ;
        RECT 4.35 0.95 4.75 1.45 ;
        RECT 2.95 1 4.75 1.3 ;
        RECT 2.95 0.95 3.45 1.35 ;
      LAYER Via1 ;
        RECT 3.07 1.02 3.33 1.28 ;
        RECT 4.42 4.27 4.68 4.53 ;
        RECT 4.42 1.07 4.68 1.33 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.5 1.95 4.15 2.2 ;
      RECT 3.9 1.05 4.15 2.2 ;
      RECT 2.2 1.05 2.45 2.2 ;
      RECT 0.5 1.05 0.75 2.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai22_1

MACRO gf180mcu_osu_sc_gp12t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai31_1 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 3.85 5.55 4.1 8.3 ;
        RECT 1.05 5.55 1.3 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 2.25 0 2.5 1.6 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.95 2.95 1.45 3.25 ;
      LAYER Metal2 ;
        RECT 0.95 2.9 1.45 3.3 ;
      LAYER Via1 ;
        RECT 1.07 2.97 1.33 3.23 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 2.95 2.3 3.25 ;
      LAYER Metal2 ;
        RECT 1.8 2.9 2.3 3.3 ;
      LAYER Via1 ;
        RECT 1.92 2.97 2.18 3.23 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.55 4.25 3.05 4.55 ;
      LAYER Metal2 ;
        RECT 2.55 4.2 3.05 4.6 ;
      LAYER Via1 ;
        RECT 2.67 4.27 2.93 4.53 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 2.95 3.6 3.25 ;
      LAYER Metal2 ;
        RECT 3.1 2.9 3.6 3.3 ;
      LAYER Via1 ;
        RECT 3.22 2.97 3.48 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 4.9 4.25 5.2 ;
        RECT 3.95 1.05 4.2 2.6 ;
        RECT 3.85 2.35 4.1 5.2 ;
        RECT 3 4.9 3.25 7.25 ;
      LAYER Metal2 ;
        RECT 3.75 4.85 4.25 5.25 ;
      LAYER Via1 ;
        RECT 3.87 4.92 4.13 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.85 3.35 2.1 ;
      RECT 3.1 1.05 3.35 2.1 ;
      RECT 1.4 1.05 1.65 2.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai31_1

MACRO gf180mcu_osu_sc_gp12t3v3__or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__or2_1 0 0 ;
  SIZE 3.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.8 8.3 ;
        RECT 1.95 5.55 2.35 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.8 0.7 ;
        RECT 2.1 0 2.35 1.9 ;
        RECT 0.4 0 0.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.9 3.6 1.4 3.9 ;
      LAYER Metal2 ;
        RECT 0.9 3.55 1.4 3.95 ;
      LAYER Via1 ;
        RECT 1.02 3.62 1.28 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.65 2.95 2.15 3.25 ;
      LAYER Metal2 ;
        RECT 1.65 2.9 2.15 3.3 ;
      LAYER Via1 ;
        RECT 1.77 2.97 2.03 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.95 4.9 3.45 5.2 ;
        RECT 2.95 1.05 3.2 7.25 ;
      LAYER Metal2 ;
        RECT 2.95 4.85 3.45 5.25 ;
      LAYER Via1 ;
        RECT 3.07 4.92 3.33 5.18 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 2.2 4.2 2.7 4.6 ;
    LAYER Via1 ;
      RECT 2.32 4.27 2.58 4.53 ;
    LAYER Metal1 ;
      RECT 0.55 5.35 0.8 7.25 ;
      RECT 0.4 2.3 0.65 5.6 ;
      RECT 0.4 4.25 2.7 4.55 ;
      RECT 0.4 2.3 1.5 2.55 ;
      RECT 1.25 1.05 1.5 2.55 ;
  END
END gf180mcu_osu_sc_gp12t3v3__or2_1

MACRO gf180mcu_osu_sc_gp12t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tbuf_1 0 0 ;
  SIZE 5.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.2 8.3 ;
        RECT 3.55 5.55 3.8 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.2 0.7 ;
        RECT 3.55 0 3.8 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 2.35 3.5 2.65 ;
      LAYER Metal2 ;
        RECT 3 2.3 3.5 2.7 ;
      LAYER Via1 ;
        RECT 3.12 2.37 3.38 2.63 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.8 5.55 3.05 7.25 ;
        RECT 1.95 1.65 3.05 1.9 ;
        RECT 2.8 1.05 3.05 1.9 ;
        RECT 2.45 3.6 2.95 3.9 ;
        RECT 1.95 4.35 2.8 4.6 ;
        RECT 2.55 2.85 2.8 4.6 ;
        RECT 1.95 5.55 3.05 5.8 ;
        RECT 1.95 2.85 2.8 3.1 ;
        RECT 1.95 4.35 2.2 5.8 ;
        RECT 1.95 1.65 2.2 3.1 ;
      LAYER Metal2 ;
        RECT 2.45 3.55 2.95 3.95 ;
      LAYER Via1 ;
        RECT 2.57 3.62 2.83 3.88 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 4.3 4.85 4.8 5.25 ;
      RECT 2.45 4.85 2.95 5.25 ;
      RECT 2.45 4.9 4.8 5.2 ;
    LAYER Via1 ;
      RECT 4.42 4.92 4.68 5.18 ;
      RECT 2.57 4.92 2.83 5.18 ;
    LAYER Metal1 ;
      RECT 4.4 1.05 4.65 7.25 ;
      RECT 4.3 4.9 4.8 5.2 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3.45 2 3.75 ;
      RECT 2.45 4.9 2.95 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tbuf_1

MACRO gf180mcu_osu_sc_gp12t3v3__tieh
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tieh 0 0 ;
  SIZE 2.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.2 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.2 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 4.9 1.8 5.2 ;
        RECT 1.4 4.85 1.65 7.25 ;
      LAYER Metal2 ;
        RECT 1.3 4.85 1.8 5.25 ;
      LAYER Via1 ;
        RECT 1.42 4.92 1.68 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.15 2.3 1.65 2.55 ;
      RECT 1.4 1.05 1.65 2.55 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tieh

MACRO gf180mcu_osu_sc_gp12t3v3__tiel
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tiel 0 0 ;
  SIZE 2.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.2 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.2 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 2.2 1.8 2.5 ;
        RECT 1.4 1.05 1.65 2.55 ;
      LAYER Metal2 ;
        RECT 1.3 2.15 1.8 2.55 ;
      LAYER Via1 ;
        RECT 1.42 2.22 1.68 2.48 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 4.95 1.65 7.25 ;
      RECT 1.15 4.95 1.65 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tiel

MACRO gf180mcu_osu_sc_gp12t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tinv_1 0 0 ;
  SIZE 3.65 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.65 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.65 0.7 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 4.9 1.95 5.2 ;
      LAYER Metal2 ;
        RECT 1.45 4.85 1.95 5.25 ;
      LAYER Via1 ;
        RECT 1.57 4.92 1.83 5.18 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.3 3.2 2.6 ;
        RECT 1 2.3 1.5 2.6 ;
      LAYER Metal2 ;
        RECT 2.7 2.25 3.2 2.65 ;
        RECT 1 2.3 3.2 2.6 ;
        RECT 1 2.25 1.5 2.65 ;
      LAYER Via1 ;
        RECT 1.12 2.32 1.38 2.58 ;
        RECT 2.82 2.32 3.08 2.58 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.8 5.55 3.05 7.25 ;
        RECT 2.2 1.65 3.05 1.9 ;
        RECT 2.8 1.05 3.05 1.9 ;
        RECT 2.2 5.55 3.05 5.8 ;
        RECT 2.05 3.6 2.6 3.9 ;
        RECT 2.2 1.65 2.45 5.8 ;
      LAYER Metal2 ;
        RECT 2.05 3.55 2.55 3.95 ;
      LAYER Via1 ;
        RECT 2.17 3.62 2.43 3.88 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 2.7 4.85 3.2 5.25 ;
      RECT 2.8 4.25 3.1 5.25 ;
      RECT 0.35 4.2 0.85 4.6 ;
      RECT 0.35 4.25 3.1 4.55 ;
    LAYER Via1 ;
      RECT 2.82 4.92 3.08 5.18 ;
      RECT 0.47 4.27 0.73 4.53 ;
    LAYER Metal1 ;
      RECT 0.55 5.55 0.8 7.25 ;
      RECT 0.5 1.9 0.75 5.8 ;
      RECT 0.35 4.25 0.85 4.55 ;
      RECT 0.55 1.05 0.8 2.15 ;
      RECT 2.7 4.9 3.2 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tinv_1

MACRO gf180mcu_osu_sc_gp12t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xnor2_1 0 0 ;
  SIZE 6.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 6.2 8.3 ;
        RECT 4.5 5.55 4.75 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 6.2 0.7 ;
        RECT 4.5 0 4.75 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 3.6 4.05 3.9 ;
        RECT 1.25 2.3 1.75 2.6 ;
      LAYER Metal2 ;
        RECT 3.6 3.55 4 3.95 ;
        RECT 3.65 1 3.95 4 ;
        RECT 1.35 1 3.95 1.3 ;
        RECT 1.3 2.25 1.7 2.65 ;
        RECT 1.35 1 1.65 2.7 ;
      LAYER Via1 ;
        RECT 1.37 2.32 1.63 2.58 ;
        RECT 3.67 3.62 3.93 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.35 2.3 4.85 2.6 ;
      LAYER Metal2 ;
        RECT 4.35 2.3 4.85 2.6 ;
        RECT 4.4 2.25 4.8 2.65 ;
        RECT 4.45 2.2 4.75 2.7 ;
      LAYER Via1 ;
        RECT 4.47 2.32 4.73 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 1.5 3.2 2.05 ;
        RECT 2.95 1.05 3.2 2.05 ;
        RECT 2.95 5.4 3.2 7.25 ;
        RECT 2.9 5.4 3.2 5.95 ;
      LAYER Metal2 ;
        RECT 2.8 1.6 3.3 2 ;
        RECT 2.85 5.5 3.25 5.9 ;
        RECT 2.9 1.6 3.2 6.05 ;
      LAYER Via1 ;
        RECT 2.92 5.57 3.18 5.83 ;
        RECT 2.92 1.67 3.18 1.93 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5.35 1.05 5.6 7.25 ;
      RECT 2.55 4.25 5.6 4.55 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3.6 3.3 3.9 ;
      RECT 3 2.3 3.3 3.9 ;
      RECT 2.9 2.3 3.4 2.6 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xnor2_1

MACRO gf180mcu_osu_sc_gp12t3v3__xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xor2_1 0 0 ;
  SIZE 6.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 6.2 8.3 ;
        RECT 4.5 5.55 4.75 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 6.2 0.7 ;
        RECT 4.5 0 4.75 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.25 2.3 1.75 2.6 ;
      LAYER Metal2 ;
        RECT 1.25 2.3 1.75 2.6 ;
        RECT 1.3 2.25 1.7 2.65 ;
      LAYER Via1 ;
        RECT 1.37 2.32 1.63 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 3.6 5.1 3.9 ;
      LAYER Metal2 ;
        RECT 4.6 3.6 5.1 3.9 ;
        RECT 4.65 3.55 5.05 3.95 ;
        RECT 1.95 3.6 2.45 3.9 ;
        RECT 2 3.55 2.4 3.95 ;
      LAYER Via1 ;
        RECT 2.07 3.62 2.33 3.88 ;
        RECT 4.72 3.62 4.98 3.88 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 1.5 3.2 2.05 ;
        RECT 2.95 1.05 3.2 2.05 ;
        RECT 2.95 5.45 3.2 7.25 ;
        RECT 2.9 5.45 3.2 5.95 ;
      LAYER Metal2 ;
        RECT 2.8 1.6 3.3 2 ;
        RECT 2.85 5.5 3.25 5.9 ;
        RECT 2.9 1.6 3.2 6.05 ;
      LAYER Via1 ;
        RECT 2.92 5.57 3.18 5.83 ;
        RECT 2.92 1.67 3.18 1.93 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5.35 1.05 5.6 7.25 ;
      RECT 2.55 4.9 5.6 5.2 ;
      RECT 4.05 2.3 5.6 2.6 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 4.25 4.05 4.55 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xor2_1

END LIBRARY
