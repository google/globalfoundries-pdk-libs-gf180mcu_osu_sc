# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_or2_1 0 0 ;
  SIZE 3.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.8 8.1 ;
        RECT 1.95 5.45 2.35 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 3.5 1.4 3.8 ;
      LAYER MET2 ;
        RECT 0.9 3.45 1.4 3.85 ;
      LAYER VIA12 ;
        RECT 1.02 3.52 1.28 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.85 2.15 3.15 ;
      LAYER MET2 ;
        RECT 1.65 2.8 2.15 3.2 ;
      LAYER VIA12 ;
        RECT 1.77 2.87 2.03 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 4.8 3.45 5.1 ;
        RECT 2.95 0.95 3.2 7.15 ;
      LAYER MET2 ;
        RECT 2.95 4.75 3.45 5.15 ;
      LAYER VIA12 ;
        RECT 3.07 4.82 3.33 5.08 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.2 4.1 2.7 4.5 ;
    LAYER VIA12 ;
      RECT 2.32 4.17 2.58 4.43 ;
    LAYER MET1 ;
      RECT 0.55 5.25 0.8 7.15 ;
      RECT 0.4 2.2 0.65 5.5 ;
      RECT 0.4 4.15 2.7 4.45 ;
      RECT 0.4 2.2 1.5 2.45 ;
      RECT 1.25 0.95 1.5 2.45 ;
  END
END gf180mcu_osu_sc_12T_or2_1
