magic
tech gf180mcuC
timestamp 1659966706
<< nwell >>
rect 0 97 88 159
<< metal1 >>
rect 0 147 88 159
rect 0 -3 88 9
<< labels >>
rlabel metal1 6 153 6 153 1 VDD
rlabel metal1 6 3 6 3 1 GND
<< end >>
