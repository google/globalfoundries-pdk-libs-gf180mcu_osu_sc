magic
tech gf180mcuC
timestamp 1659987912
<< nwell >>
rect -17 97 44 159
<< nmos >>
rect 2 16 8 33
rect 19 16 25 33
<< pmos >>
rect 2 106 8 140
rect 19 106 25 140
<< ndiff >>
rect -8 31 2 33
rect -8 18 -6 31
rect -1 18 2 31
rect -8 16 2 18
rect 8 31 19 33
rect 8 18 11 31
rect 16 18 19 31
rect 8 16 19 18
rect 25 31 35 33
rect 25 18 28 31
rect 33 18 35 31
rect 25 16 35 18
<< pdiff >>
rect -8 138 2 140
rect -8 108 -6 138
rect -1 108 2 138
rect -8 106 2 108
rect 8 138 19 140
rect 8 108 11 138
rect 16 108 19 138
rect 8 106 19 108
rect 25 138 35 140
rect 25 108 28 138
rect 33 108 35 138
rect 25 106 35 108
<< ndiffc >>
rect -6 18 -1 31
rect 11 18 16 31
rect 28 18 33 31
<< pdiffc >>
rect -6 108 -1 138
rect 11 108 16 138
rect 28 108 33 138
<< psubdiff >>
rect -8 7 2 9
rect -8 2 -6 7
rect -1 2 2 7
rect -8 0 2 2
rect 16 7 26 9
rect 16 2 18 7
rect 23 2 26 7
rect 16 0 26 2
<< nsubdiff >>
rect -8 154 2 156
rect -8 149 -6 154
rect -1 149 2 154
rect -8 147 2 149
rect 16 154 26 156
rect 16 149 18 154
rect 23 149 26 154
rect 16 147 26 149
<< psubdiffcont >>
rect -6 2 -1 7
rect 18 2 23 7
<< nsubdiffcont >>
rect -6 149 -1 154
rect 18 149 23 154
<< polysilicon >>
rect 2 140 8 145
rect 19 140 25 145
rect 2 88 8 106
rect 2 86 14 88
rect 2 80 6 86
rect 12 80 14 86
rect 2 78 14 80
rect 2 33 8 78
rect 19 64 25 106
rect 13 61 25 64
rect 13 55 15 61
rect 21 55 25 61
rect 13 52 25 55
rect 19 33 25 52
rect 2 11 8 16
rect 19 11 25 16
<< polycontact >>
rect 6 80 12 86
rect 15 55 21 61
<< metal1 >>
rect -17 154 44 159
rect -17 148 -6 154
rect 0 148 18 154
rect 24 148 44 154
rect -17 147 44 148
rect -6 138 -1 140
rect -6 61 -1 108
rect 11 138 16 147
rect 11 106 16 108
rect 28 138 33 140
rect 28 99 33 108
rect 26 93 28 99
rect 34 93 36 99
rect 4 80 6 86
rect 12 80 14 86
rect -6 55 15 61
rect 21 55 23 61
rect -6 31 -1 55
rect -6 16 -1 18
rect 11 31 16 33
rect 11 9 16 18
rect 28 31 33 93
rect 28 16 33 18
rect -17 8 44 9
rect -17 2 -6 8
rect 0 2 18 8
rect 24 2 44 8
rect -17 -3 44 2
<< via1 >>
rect -6 149 -1 154
rect -1 149 0 154
rect -6 148 0 149
rect 18 149 23 154
rect 23 149 24 154
rect 18 148 24 149
rect 28 93 34 99
rect 6 80 12 86
rect -6 7 0 8
rect -6 2 -1 7
rect -1 2 0 7
rect 18 7 24 8
rect 18 2 23 7
rect 23 2 24 7
<< metal2 >>
rect -7 154 1 155
rect 17 154 25 155
rect -8 148 -6 154
rect 0 148 2 154
rect 16 148 18 154
rect 24 148 26 154
rect -7 147 1 148
rect 17 147 25 148
rect 26 99 36 100
rect 26 93 28 99
rect 34 93 36 99
rect 26 92 36 93
rect 5 86 13 87
rect 4 80 6 86
rect 12 80 14 86
rect 5 79 13 80
rect -7 8 1 9
rect 17 8 25 9
rect -8 2 -6 8
rect 0 2 2 8
rect 16 2 18 8
rect 24 2 26 8
rect -7 1 1 2
rect 17 1 25 2
<< labels >>
rlabel metal2 -3 5 -3 5 1 GND
rlabel metal2 -3 151 -3 151 1 VDD
rlabel metal2 31 96 31 96 1 Y
port 2 n
rlabel metal2 9 83 9 83 1 A
port 1 n
<< end >>
