# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__oai22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai22_1 0 0 ;
  SIZE 5.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.5 6.15 ;
        RECT 3.6 3.5 3.85 6.15 ;
        RECT 0.65 3.5 0.9 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.5 0.6 ;
        RECT 1.35 0 1.6 1.45 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 2.2 1.2 2.5 ;
      LAYER MET2 ;
        RECT 0.7 2.15 1.2 2.55 ;
      LAYER VIA12 ;
        RECT 0.82 2.22 1.08 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.2 2.15 2.5 ;
      LAYER MET2 ;
        RECT 1.65 2.15 2.15 2.55 ;
      LAYER VIA12 ;
        RECT 1.77 2.22 2.03 2.48 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 2.2 3.05 2.5 ;
      LAYER MET2 ;
        RECT 2.55 2.15 3.05 2.55 ;
      LAYER VIA12 ;
        RECT 2.67 2.22 2.93 2.48 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 2.2 3.85 2.5 ;
      LAYER MET2 ;
        RECT 3.35 2.15 3.85 2.55 ;
      LAYER VIA12 ;
        RECT 3.47 2.22 3.73 2.48 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.5 0.85 5 1.15 ;
        RECT 2.1 2.75 4.9 3.05 ;
        RECT 4.6 0.85 4.9 3.05 ;
        RECT 2.1 2.75 2.45 5.2 ;
        RECT 3.05 0.85 3.55 1.2 ;
        RECT 3.15 0.85 3.4 1.45 ;
      LAYER MET2 ;
        RECT 3.05 0.85 5 1.15 ;
        RECT 4.55 0.8 4.95 1.2 ;
        RECT 3.05 0.8 3.55 1.2 ;
      LAYER VIA12 ;
        RECT 3.17 0.87 3.43 1.13 ;
        RECT 4.62 0.87 4.88 1.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.7 4.25 1.95 ;
      RECT 4 0.95 4.25 1.95 ;
      RECT 2.2 0.95 2.55 1.95 ;
      RECT 0.5 0.95 0.75 1.95 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai22_1
