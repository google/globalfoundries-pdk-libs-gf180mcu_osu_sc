# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_clkbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_clkbuf_4 0 0 ;
  SIZE 5.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.6 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.6 0.6 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 4.85 4.35 5.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 2.05 4.2 2.3 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 3.85 4.8 4.35 5.2 ;
        RECT 3.8 4.85 4.35 5.15 ;
      LAYER VIA12 ;
        RECT 3.97 4.87 4.23 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_12T_clkbuf_4
