# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_8 0 0 ;
  SIZE 11.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 11.5 6.15 ;
        RECT 10.7 3.5 10.95 6.15 ;
        RECT 8.95 3.5 9.2 6.15 ;
        RECT 7.25 3.5 7.5 6.15 ;
        RECT 5.55 3.5 5.8 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 1.1 3.5 1.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 11.5 0.6 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.95 0 9.2 1.8 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.1 0 1.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 1.45 2.25 2.9 ;
      LAYER MET2 ;
        RECT 1.85 1.5 2.35 1.9 ;
      LAYER VIA12 ;
        RECT 1.97 1.57 2.23 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.8 3.5 10.45 3.8 ;
        RECT 9.8 0.95 10.05 5.2 ;
        RECT 4.7 3 10.05 3.25 ;
        RECT 4.7 2.05 10.05 2.3 ;
        RECT 8.1 0.95 8.35 5.2 ;
        RECT 6.4 0.95 6.65 5.2 ;
        RECT 4.7 0.95 4.95 5.2 ;
      LAYER MET2 ;
        RECT 9.95 3.5 10.45 3.8 ;
        RECT 10 3.45 10.4 3.85 ;
      LAYER VIA12 ;
        RECT 10.07 3.52 10.33 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.4 2.8 3.95 3.2 ;
    LAYER VIA12 ;
      RECT 3.57 2.87 3.83 3.13 ;
      RECT 2.52 2.87 2.78 3.13 ;
    LAYER MET1 ;
      RECT 3 3.5 3.25 5.2 ;
      RECT 3.05 2.2 3.3 3.7 ;
      RECT 4.15 2.1 4.4 2.55 ;
      RECT 3 0.95 3.25 2.55 ;
      RECT 3 2.2 4.4 2.45 ;
      RECT 2.5 0.95 2.75 5.2 ;
      RECT 2.5 2.75 2.8 3.25 ;
      RECT 3.55 2.75 3.85 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_8
