*
* Filename: test.sp
* Author: James E. Stine, Jr.
* Course: none
* Credits: none
* Title: GF180 MCU inverter test

***********************************************************************
* Parameters and models
***********************************************************************
.inc "/home/jstine/Desktop/gf180/mcu/018MCU/MODEL/Hspice/YI-141-SM064/Rev9/design.hspice"
.lib "/home/jstine/Desktop/gf180/mcu/018MCU/MODEL/Hspice/YI-141-SM064/Rev9/sm141064.hspice" typical
.temp 25
.param SUPPLY=3.3V

***********************************************************************
* Simulation netlist
***********************************************************************
Vdd	vdd	gnd	'SUPPLY'
Vin	A	gnd	PULSE	0 'SUPPLY' 0ps 25p 25p 500p 1000p

.option scale=0.05u
.subckt gf180mcu_osu_sc_12T_inv_1 A Y
X0 Y A VDD VDD pmos_3p3 w=34 l=6
X1 Y A GND GND nmos_3p3 w=17 l=6
.ends

***********************************************************************
* Stimulus
***********************************************************************

.dc Vin 0V +5V 100mV
.tran .05n 5n 

.probe v(A) v(Out)
.op
.options probe post acct list node measout captab
.end
