# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_tinv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_tinv_2 0 0 ;
  SIZE 6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 6 8.1 ;
        RECT 5.05 5.45 5.3 8.1 ;
        RECT 3.3 5.45 3.55 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6 0.6 ;
        RECT 5 0 5.25 1.8 ;
        RECT 3.3 0 3.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 3.5 1.45 3.8 ;
      LAYER MET2 ;
        RECT 0.95 3.45 1.45 3.85 ;
      LAYER VIA12 ;
        RECT 1.07 3.52 1.33 3.78 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 2.2 1.25 2.5 ;
      LAYER MET2 ;
        RECT 0.75 2.15 1.25 2.55 ;
      LAYER VIA12 ;
        RECT 0.87 2.22 1.13 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 4.8 1.25 5.1 ;
      LAYER MET2 ;
        RECT 0.75 4.75 1.25 5.15 ;
      LAYER VIA12 ;
        RECT 0.87 4.82 1.13 5.08 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.15 4.15 4.75 4.45 ;
        RECT 4.15 4 4.6 4.55 ;
        RECT 4.15 0.95 4.4 7.15 ;
      LAYER MET2 ;
        RECT 4.25 4.1 4.75 4.5 ;
      LAYER VIA12 ;
        RECT 4.37 4.17 4.63 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 1.8 4.75 3.35 5.15 ;
    LAYER VIA12 ;
      RECT 2.97 4.82 3.23 5.08 ;
      RECT 1.92 4.82 2.18 5.08 ;
    LAYER MET1 ;
      RECT 2.45 0.95 2.7 7.15 ;
      RECT 3.6 3.45 3.85 3.9 ;
      RECT 2.45 3.55 3.85 3.85 ;
      RECT 1.95 0.95 2.2 7.15 ;
      RECT 1.9 4.7 2.2 5.2 ;
      RECT 2.95 4.7 3.25 5.2 ;
  END
END gf180mcu_osu_sc_12T_tinv_2
