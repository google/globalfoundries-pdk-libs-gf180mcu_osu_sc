# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dlat_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dlat_1 0 0 ;
  SIZE 9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal2 ;
        RECT 5.2 4.2 5.7 4.6 ;
        RECT 3.45 4.25 5.7 4.55 ;
        RECT 3.5 4.2 3.9 4.6 ;
      LAYER Metal1 ;
        RECT 5.2 4.25 5.7 4.55 ;
        RECT 3.45 4.25 3.95 4.55 ;
      LAYER Via1 ;
        RECT 3.57 4.27 3.83 4.53 ;
        RECT 5.32 4.27 5.58 4.53 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 9 8.3 ;
        RECT 7.3 5.55 7.55 8.3 ;
        RECT 4.85 5.55 5.1 8.3 ;
        RECT 1.45 6.35 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 9 0.7 ;
        RECT 7.3 0 7.55 1.9 ;
        RECT 4.7 0 5.1 1.9 ;
        RECT 1.45 0 1.85 1.9 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1.85 4.2 2.35 4.6 ;
      LAYER Metal1 ;
        RECT 1.85 4.25 2.35 4.55 ;
      LAYER Via1 ;
        RECT 1.97 4.27 2.23 4.53 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 8.15 4.9 8.65 5.2 ;
        RECT 8.2 4.85 8.6 5.25 ;
      LAYER Metal1 ;
        RECT 8.15 4.9 8.65 5.2 ;
        RECT 8.15 4.85 8.55 5.25 ;
        RECT 8.15 1.05 8.4 7.25 ;
      LAYER Via1 ;
        RECT 8.27 4.92 8.53 5.18 ;
    END
  END Q
  OBS
    LAYER Metal2 ;
      RECT 6.75 3.55 7.25 3.95 ;
      RECT 4.55 3.55 4.95 3.95 ;
      RECT 0.35 3.55 0.85 3.95 ;
      RECT 0.35 3.6 7.25 3.9 ;
      RECT 6.5 4.85 6.9 5.25 ;
      RECT 6.45 4.9 6.95 5.2 ;
    LAYER Via1 ;
      RECT 6.87 3.62 7.13 3.88 ;
      RECT 6.57 4.92 6.83 5.18 ;
      RECT 4.62 3.62 4.88 3.88 ;
      RECT 0.47 3.62 0.73 3.88 ;
    LAYER Metal1 ;
      RECT 6.45 4.85 6.7 7.25 ;
      RECT 6.45 4.85 6.85 5.4 ;
      RECT 6.45 4.9 6.95 5.2 ;
      RECT 6.45 4.9 7.8 5.15 ;
      RECT 7.5 2.15 7.8 5.15 ;
      RECT 6.45 2.15 7.8 2.4 ;
      RECT 6.45 1.05 6.7 2.4 ;
      RECT 5.7 5.35 5.95 7.25 ;
      RECT 5.95 2.05 6.2 5.6 ;
      RECT 2.6 4.8 3.1 5.1 ;
      RECT 2.7 2.65 3 5.1 ;
      RECT 2.7 2.65 6.2 2.95 ;
      RECT 5.7 1.05 5.95 2.3 ;
      RECT 3.15 5.55 3.4 7.25 ;
      RECT 1.15 5.55 3.4 5.8 ;
      RECT 1.15 2.15 1.4 5.8 ;
      RECT 1.1 4.25 1.55 4.55 ;
      RECT 1.15 2.15 3.4 2.4 ;
      RECT 3.15 1.05 3.4 2.4 ;
      RECT 0.6 1.05 0.85 7.25 ;
      RECT 0.5 3.55 0.85 3.95 ;
      RECT 0.35 3.6 0.85 3.9 ;
      RECT 0.45 3.55 0.85 3.9 ;
      RECT 6.75 3.6 7.25 3.9 ;
      RECT 4.5 3.6 5 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dlat_1
