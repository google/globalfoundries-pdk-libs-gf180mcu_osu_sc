magic
tech gf180mcuC
timestamp 1661875450
<< nwell >>
rect 0 61 44 123
<< nmos >>
rect 19 19 25 36
<< pmos >>
rect 19 70 25 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 35 36
rect 25 21 28 34
rect 33 21 35 34
rect 25 19 35 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 35 104
rect 25 77 28 102
rect 33 77 35 102
rect 25 70 35 77
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
<< pdiffc >>
rect 11 72 16 102
rect 28 77 33 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
<< psubdiffcont >>
rect 11 5 16 10
<< nsubdiffcont >>
rect 11 113 16 118
<< polysilicon >>
rect 19 104 25 109
rect 19 51 25 70
rect 19 49 33 51
rect 19 44 26 49
rect 31 44 33 49
rect 19 42 33 44
rect 19 36 25 42
rect 19 14 25 19
<< polycontact >>
rect 26 44 31 49
<< metal1 >>
rect 0 118 44 123
rect 0 112 11 118
rect 17 112 44 118
rect 0 111 44 112
rect 11 102 16 111
rect 28 102 33 104
rect 28 76 33 77
rect 11 70 16 72
rect 26 70 28 76
rect 34 70 36 76
rect 28 69 33 70
rect 23 44 26 49
rect 31 44 33 49
rect 11 34 16 36
rect 11 12 16 21
rect 28 34 33 44
rect 28 19 33 21
rect 0 11 44 12
rect 0 5 11 11
rect 17 5 44 11
rect 0 0 44 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 28 70 34 76
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
<< metal2 >>
rect 10 118 18 119
rect 9 112 11 118
rect 17 112 19 118
rect 10 111 18 112
rect 26 76 36 77
rect 26 70 28 76
rect 34 70 36 76
rect 26 69 36 70
rect 10 11 18 12
rect 9 5 11 11
rect 17 5 19 11
rect 10 4 18 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 31 73 31 73 1 Y
port 2 n
<< end >>
