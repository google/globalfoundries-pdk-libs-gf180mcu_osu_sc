# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_aoi22_1 0 0 ;
  SIZE 5.4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.4 6.15 ;
        RECT 1.4 4.25 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.4 0.6 ;
        RECT 3.5 0 3.75 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.4 2.85 2.9 3.15 ;
      LAYER MET2 ;
        RECT 2.4 2.8 2.9 3.2 ;
      LAYER VIA12 ;
        RECT 2.52 2.87 2.78 3.13 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 2.85 3.8 3.15 ;
      LAYER MET2 ;
        RECT 3.3 2.8 3.8 3.2 ;
      LAYER VIA12 ;
        RECT 3.42 2.87 3.68 3.13 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.5 4.05 4.8 4.55 ;
        RECT 4.55 2.05 4.8 4.55 ;
        RECT 2.1 2.05 4.8 2.3 ;
        RECT 2.1 0.95 2.35 2.3 ;
        RECT 3 4.15 3.5 4.45 ;
        RECT 3.1 4.15 3.35 5.2 ;
      LAYER MET2 ;
        RECT 4.45 4.05 4.85 4.55 ;
        RECT 3 4.15 4.85 4.45 ;
        RECT 3 4.1 3.5 4.5 ;
      LAYER VIA12 ;
        RECT 3.12 4.17 3.38 4.43 ;
        RECT 4.52 4.17 4.78 4.43 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.95 3.65 4.25 5.2 ;
      RECT 2.25 3.65 2.5 5.2 ;
      RECT 0.55 3.65 0.8 5.2 ;
      RECT 0.55 3.65 4.25 3.9 ;
  END
END gf180mcu_osu_sc_9T_aoi22_1
