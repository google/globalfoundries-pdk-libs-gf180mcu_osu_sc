magic
tech gf180mcuC
timestamp 1661533308
<< nwell >>
rect 0 97 134 159
<< nmos >>
rect 19 55 25 72
rect 36 55 42 72
rect 52 55 58 72
rect 75 55 81 72
rect 91 55 97 72
rect 108 55 114 72
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 52 106 58 140
rect 75 106 81 140
rect 91 106 97 140
rect 108 106 114 140
<< ndiff >>
rect 9 70 19 72
rect 9 57 11 70
rect 16 57 19 70
rect 9 55 19 57
rect 25 70 36 72
rect 25 57 28 70
rect 33 57 36 70
rect 25 55 36 57
rect 42 55 52 72
rect 58 62 75 72
rect 58 57 64 62
rect 69 57 75 62
rect 58 55 75 57
rect 81 55 91 72
rect 97 69 108 72
rect 97 57 100 69
rect 105 57 108 69
rect 97 55 108 57
rect 114 70 124 72
rect 114 57 117 70
rect 122 57 124 70
rect 114 55 124 57
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 114 28 138
rect 33 114 36 138
rect 25 106 36 114
rect 42 106 52 140
rect 58 138 75 140
rect 58 133 64 138
rect 69 133 75 138
rect 58 106 75 133
rect 81 106 91 140
rect 97 138 108 140
rect 97 114 100 138
rect 105 114 108 138
rect 97 106 108 114
rect 114 138 124 140
rect 114 108 117 138
rect 122 108 124 138
rect 114 106 124 108
<< ndiffc >>
rect 11 57 16 70
rect 28 57 33 70
rect 64 57 69 62
rect 100 57 105 69
rect 117 57 122 70
<< pdiffc >>
rect 11 108 16 138
rect 28 114 33 138
rect 64 133 69 138
rect 100 114 105 138
rect 117 108 122 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
rect 57 46 66 48
rect 57 41 59 46
rect 64 41 66 46
rect 57 39 66 41
rect 81 46 90 48
rect 81 41 83 46
rect 88 41 90 46
rect 81 39 90 41
rect 105 46 114 48
rect 105 41 107 46
rect 112 41 114 46
rect 105 39 114 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
rect 81 154 90 156
rect 81 149 83 154
rect 88 149 90 154
rect 81 147 90 149
rect 105 154 114 156
rect 105 149 107 154
rect 112 149 114 154
rect 105 147 114 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
rect 59 41 64 46
rect 83 41 88 46
rect 107 41 112 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
rect 83 149 88 154
rect 107 149 112 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 52 140 58 145
rect 75 140 81 145
rect 91 140 97 145
rect 108 140 114 145
rect 19 104 25 106
rect 36 104 42 106
rect 19 99 42 104
rect 52 104 58 106
rect 75 104 81 106
rect 52 102 62 104
rect 19 88 25 99
rect 52 97 54 102
rect 60 97 62 102
rect 52 95 62 97
rect 71 102 81 104
rect 71 96 73 102
rect 79 96 81 102
rect 91 104 97 106
rect 108 104 114 106
rect 91 99 114 104
rect 71 94 81 96
rect 19 86 32 88
rect 19 80 24 86
rect 30 80 32 86
rect 19 78 32 80
rect 47 82 58 84
rect 19 74 42 78
rect 47 76 49 82
rect 55 76 58 82
rect 47 74 58 76
rect 19 72 25 74
rect 36 72 42 74
rect 52 72 58 74
rect 75 72 81 94
rect 87 92 97 94
rect 87 87 89 92
rect 95 87 97 92
rect 108 88 114 99
rect 87 85 97 87
rect 91 72 97 85
rect 102 86 114 88
rect 102 80 104 86
rect 110 80 114 86
rect 102 78 114 80
rect 108 72 114 78
rect 19 50 25 55
rect 36 50 42 55
rect 52 50 58 55
rect 75 50 81 55
rect 91 50 97 55
rect 108 50 114 55
<< polycontact >>
rect 54 97 60 102
rect 73 96 79 102
rect 24 80 30 86
rect 49 76 55 82
rect 89 87 95 92
rect 104 80 110 86
<< metal1 >>
rect 0 154 134 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 83 154
rect 89 148 107 154
rect 113 148 134 154
rect 0 147 134 148
rect 11 138 16 140
rect 28 138 33 147
rect 64 138 69 140
rect 64 127 69 133
rect 63 125 69 127
rect 100 138 105 147
rect 61 119 63 125
rect 69 119 71 125
rect 28 112 33 114
rect 11 101 16 108
rect 54 109 94 114
rect 100 112 105 114
rect 117 138 122 140
rect 54 102 60 109
rect 89 104 94 109
rect 117 104 122 108
rect 73 102 79 104
rect 11 96 47 101
rect 52 97 54 102
rect 60 97 62 102
rect 11 70 16 96
rect 41 92 47 96
rect 73 92 79 96
rect 89 98 122 104
rect 89 93 95 98
rect 41 87 79 92
rect 87 92 97 93
rect 87 87 89 92
rect 95 87 97 92
rect 22 80 24 86
rect 30 80 32 86
rect 102 82 104 86
rect 47 76 49 82
rect 55 80 104 82
rect 110 80 112 86
rect 55 76 109 80
rect 11 55 16 57
rect 28 70 33 72
rect 63 70 69 71
rect 61 64 63 70
rect 69 64 71 70
rect 100 69 105 71
rect 63 62 69 64
rect 28 48 33 57
rect 64 55 69 57
rect 100 48 105 57
rect 117 70 122 98
rect 117 55 122 57
rect 0 47 134 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 59 47
rect 65 41 83 47
rect 89 41 107 47
rect 113 41 134 47
rect 0 36 134 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 83 149 88 154
rect 88 149 89 154
rect 83 148 89 149
rect 107 149 112 154
rect 112 149 113 154
rect 107 148 113 149
rect 63 119 69 125
rect 24 80 30 86
rect 104 80 110 86
rect 63 64 69 70
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
rect 59 46 65 47
rect 59 41 64 46
rect 64 41 65 46
rect 83 46 89 47
rect 83 41 88 46
rect 88 41 89 46
rect 107 46 113 47
rect 107 41 112 46
rect 112 41 113 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 81 148 83 154
rect 89 148 91 154
rect 105 148 107 154
rect 113 148 115 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 63 126 69 127
rect 62 125 70 126
rect 62 119 63 125
rect 69 119 70 125
rect 62 118 70 119
rect 23 86 31 87
rect 22 80 24 86
rect 30 80 32 86
rect 23 79 31 80
rect 63 71 69 118
rect 103 86 111 87
rect 102 80 104 86
rect 110 80 112 86
rect 103 79 111 80
rect 61 70 71 71
rect 61 64 63 70
rect 69 64 71 70
rect 61 63 71 64
rect 10 47 18 48
rect 34 47 42 48
rect 58 47 66 48
rect 82 47 90 48
rect 106 47 114 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 57 41 59 47
rect 65 41 67 47
rect 81 41 83 47
rect 89 41 91 47
rect 105 41 107 47
rect 113 41 115 47
rect 10 40 18 41
rect 34 40 42 41
rect 58 40 66 41
rect 82 40 90 41
rect 106 40 114 41
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 14 44 14 44 1 GND
rlabel metal2 66 121 66 121 1 Y
port 3 n
rlabel metal2 27 83 27 83 1 A
port 1 n
rlabel metal2 107 83 107 83 1 B
port 4 n
<< end >>
