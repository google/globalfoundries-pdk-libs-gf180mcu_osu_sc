* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__tbuf_8 A Y EN EN_BAR
X0 VSS a_13_19 Y VSS nmos_3p3 w=17 l=6
X1 VSS a_13_19 Y VSS nmos_3p3 w=17 l=6
X2 VSS a_13_19 Y VSS nmos_3p3 w=17 l=6
X3 Y a_13_19 VSS VSS nmos_3p3 w=17 l=6
X4 VDD a_13_19 Y VDD pmos_3p3 w=34 l=6
X5 Y a_13_19 VDD VDD pmos_3p3 w=34 l=6
X6 VDD a_13_19 Y VDD pmos_3p3 w=34 l=6
X7 VDD a_13_19 Y VDD pmos_3p3 w=34 l=6
X8 Y a_13_19 VDD VDD pmos_3p3 w=34 l=6
X9 Y a_13_19 VDD VDD pmos_3p3 w=34 l=6
X10 a_29_19 EN a_13_19 VSS nmos_3p3 w=17 l=6
X11 Y a_13_19 VSS VSS nmos_3p3 w=17 l=6
X12 Y a_13_19 VSS VSS nmos_3p3 w=17 l=6
X13 Y a_13_19 VDD VDD pmos_3p3 w=34 l=6
X14 VDD a_13_19 Y VDD pmos_3p3 w=34 l=6
X15 VDD A a_29_109 VDD pmos_3p3 w=34 l=6
X16 Y a_13_19 VSS VSS nmos_3p3 w=17 l=6
X17 VSS A a_29_19 VSS nmos_3p3 w=17 l=6
X18 VSS a_13_19 Y VSS nmos_3p3 w=17 l=6
X19 a_29_109 EN_BAR a_13_19 VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
