magic
tech gf180mcuC
timestamp 1659735289
<< nwell >>
rect 0 97 123 159
<< nmos >>
rect 19 16 25 33
rect 36 16 42 33
rect 47 16 53 33
rect 70 16 76 33
rect 81 16 87 33
rect 98 16 104 33
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 47 106 53 140
rect 70 106 76 140
rect 81 106 87 140
rect 98 106 104 140
<< ndiff >>
rect 56 33 66 34
rect 9 31 19 33
rect 9 18 11 31
rect 16 18 19 31
rect 9 16 19 18
rect 25 31 36 33
rect 25 18 28 31
rect 33 18 36 31
rect 25 16 36 18
rect 42 16 47 33
rect 53 32 70 33
rect 53 18 59 32
rect 64 18 70 32
rect 53 16 70 18
rect 76 16 81 33
rect 87 31 98 33
rect 87 18 90 31
rect 95 18 98 31
rect 87 16 98 18
rect 104 31 114 33
rect 104 18 107 31
rect 112 18 114 31
rect 104 16 114 18
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 108 28 138
rect 33 108 36 138
rect 25 106 36 108
rect 42 106 47 140
rect 53 138 70 140
rect 53 108 59 138
rect 64 108 70 138
rect 53 106 70 108
rect 76 106 81 140
rect 87 138 98 140
rect 87 108 90 138
rect 95 108 98 138
rect 87 106 98 108
rect 104 138 114 140
rect 104 108 107 138
rect 112 108 114 138
rect 104 106 114 108
<< ndiffc >>
rect 11 18 16 31
rect 28 18 33 31
rect 59 18 64 32
rect 90 18 95 31
rect 107 18 112 31
<< pdiffc >>
rect 11 108 16 138
rect 28 108 33 138
rect 59 108 64 138
rect 90 108 95 138
rect 107 108 112 138
<< psubdiff >>
rect 9 7 18 9
rect 9 2 11 7
rect 16 2 18 7
rect 9 0 18 2
rect 33 7 42 9
rect 33 2 35 7
rect 40 2 42 7
rect 33 0 42 2
rect 57 7 66 9
rect 57 2 59 7
rect 64 2 66 7
rect 57 0 66 2
rect 81 7 90 9
rect 81 2 83 7
rect 88 2 90 7
rect 81 0 90 2
rect 105 7 114 9
rect 105 2 107 7
rect 112 2 114 7
rect 105 0 114 2
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
rect 81 154 90 156
rect 81 149 83 154
rect 88 149 90 154
rect 81 147 90 149
rect 105 154 114 156
rect 105 149 107 154
rect 112 149 114 154
rect 105 147 114 149
<< psubdiffcont >>
rect 11 2 16 7
rect 35 2 40 7
rect 59 2 64 7
rect 83 2 88 7
rect 107 2 112 7
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
rect 83 149 88 154
rect 107 149 112 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 47 140 53 145
rect 70 140 76 145
rect 81 140 87 145
rect 98 140 104 145
rect 19 103 25 106
rect 36 103 42 106
rect 19 98 42 103
rect 47 101 53 106
rect 47 99 61 101
rect 19 49 25 98
rect 47 93 53 99
rect 59 93 61 99
rect 47 91 61 93
rect 70 88 76 106
rect 81 101 87 106
rect 98 101 104 106
rect 81 95 104 101
rect 69 86 81 88
rect 69 80 72 86
rect 78 80 81 86
rect 69 78 81 80
rect 39 73 53 75
rect 39 67 41 73
rect 47 67 53 73
rect 39 64 53 67
rect 47 49 53 64
rect 70 49 76 78
rect 98 75 104 95
rect 92 73 104 75
rect 92 67 94 73
rect 100 67 104 73
rect 92 65 104 67
rect 19 47 91 49
rect 19 41 27 47
rect 33 41 83 47
rect 89 41 91 47
rect 19 38 42 41
rect 19 33 25 38
rect 36 33 42 38
rect 47 33 53 41
rect 70 33 76 41
rect 81 39 91 41
rect 81 33 87 39
rect 98 33 104 65
rect 19 11 25 16
rect 36 11 42 16
rect 47 11 53 16
rect 70 11 76 16
rect 81 11 87 16
rect 98 11 104 16
<< polycontact >>
rect 53 93 59 99
rect 72 80 78 86
rect 41 67 47 73
rect 94 67 100 73
rect 27 41 33 47
rect 83 41 89 47
<< metal1 >>
rect 0 154 123 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 83 154
rect 89 148 107 154
rect 113 148 123 154
rect 0 147 123 148
rect 11 138 16 140
rect 11 86 16 108
rect 28 138 33 147
rect 59 138 64 140
rect 28 106 33 108
rect 58 112 59 114
rect 90 138 95 147
rect 90 106 95 108
rect 107 138 112 140
rect 58 104 64 106
rect 107 99 112 108
rect 51 93 53 99
rect 59 93 112 99
rect 11 80 72 86
rect 78 80 81 86
rect 11 31 16 80
rect 39 67 41 73
rect 47 67 94 73
rect 100 67 102 73
rect 107 47 112 93
rect 25 41 27 47
rect 33 41 35 47
rect 81 41 83 47
rect 89 41 112 47
rect 58 34 64 36
rect 11 16 16 18
rect 28 31 33 33
rect 58 25 59 28
rect 28 9 33 18
rect 59 16 64 18
rect 90 31 95 33
rect 90 9 95 18
rect 107 31 112 41
rect 107 16 112 18
rect 0 8 123 9
rect 0 2 11 8
rect 17 2 35 8
rect 41 2 59 8
rect 65 2 83 8
rect 89 2 107 8
rect 113 2 123 8
rect 0 -3 123 2
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 83 149 88 154
rect 88 149 89 154
rect 83 148 89 149
rect 107 149 112 154
rect 112 149 113 154
rect 107 148 113 149
rect 58 108 59 112
rect 59 108 64 112
rect 58 106 64 108
rect 41 67 47 73
rect 94 67 100 73
rect 27 41 33 47
rect 58 32 64 34
rect 58 28 59 32
rect 59 28 64 32
rect 11 7 17 8
rect 11 2 16 7
rect 16 2 17 7
rect 35 7 41 8
rect 35 2 40 7
rect 40 2 41 7
rect 59 7 65 8
rect 59 2 64 7
rect 64 2 65 7
rect 83 7 89 8
rect 83 2 88 7
rect 88 2 89 7
rect 107 7 113 8
rect 107 2 112 7
rect 112 2 113 7
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 81 148 83 154
rect 89 148 91 154
rect 105 148 107 154
rect 113 148 115 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 58 113 64 116
rect 57 112 65 113
rect 57 106 58 112
rect 64 106 65 112
rect 57 105 65 106
rect 40 73 48 74
rect 39 67 41 73
rect 47 67 49 73
rect 40 66 48 67
rect 26 47 34 48
rect 25 41 27 47
rect 33 41 35 47
rect 26 40 34 41
rect 58 35 64 105
rect 93 73 101 74
rect 92 67 94 73
rect 100 67 102 73
rect 93 66 101 67
rect 56 34 66 35
rect 56 28 58 34
rect 64 28 66 34
rect 56 27 66 28
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 82 8 90 9
rect 106 8 114 9
rect 9 2 11 8
rect 17 2 19 8
rect 33 2 35 8
rect 41 2 43 8
rect 57 2 59 8
rect 65 2 67 8
rect 81 2 83 8
rect 89 2 91 8
rect 105 2 107 8
rect 113 2 115 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
rect 82 1 90 2
rect 106 1 114 2
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 14 5 14 5 1 GND
rlabel metal2 61 108 61 108 1 Y
port 3 n
rlabel metal2 30 44 30 44 1 A
port 1 n
rlabel metal2 97 70 97 70 1 B
port 4 n
<< end >>
