# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__lshifup 0 0 ;
  SIZE 7.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 1.9 6.15 ;
        RECT 0.55 3.5 0.85 6.15 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.15 5.55 7.1 6.15 ;
        RECT 5.35 3.5 5.65 6.15 ;
        RECT 3.3 4.05 3.8 6.15 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 7.1 0.6 ;
        RECT 5.35 0 5.65 1.8 ;
        RECT 3.3 0 3.8 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.65 2.05 3.15 2.35 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 2.65 2.05 3.15 2.35 ;
        RECT 2.65 2 3.1 2.4 ;
        RECT 2.8 1.4 3.1 2.4 ;
        RECT 0.7 1.4 3.1 1.7 ;
        RECT 0.55 2.15 1.05 2.55 ;
        RECT 0.7 1.4 1 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
        RECT 2.77 2.07 3.03 2.33 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.2 2.2 6.6 2.5 ;
        RECT 6.25 0.95 6.55 5.2 ;
      LAYER MET2 ;
        RECT 6.15 2.15 6.65 2.55 ;
      LAYER VIA12 ;
        RECT 6.27 2.22 6.53 2.48 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.2 3.5 2.7 3.9 ;
      RECT 2.2 3.5 4.45 3.85 ;
      RECT 4.15 2.8 4.45 3.85 ;
      RECT 5.4 2.8 5.9 3.2 ;
      RECT 4.1 2.8 4.5 3.2 ;
      RECT 4.05 2.85 5.9 3.15 ;
      RECT 4.05 2.8 4.55 3.15 ;
      RECT 1.45 2.85 3.75 3.15 ;
      RECT 3.45 2.05 3.75 3.15 ;
      RECT 1.45 2.15 1.75 3.15 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 3.45 2.05 4.45 2.4 ;
      RECT 3.95 2 4.45 2.4 ;
    LAYER VIA12 ;
      RECT 5.52 2.87 5.78 3.13 ;
      RECT 4.17 2.87 4.43 3.13 ;
      RECT 4.07 2.07 4.33 2.33 ;
      RECT 2.32 3.57 2.58 3.83 ;
      RECT 1.47 2.22 1.73 2.48 ;
    LAYER MET1 ;
      RECT 4.4 3.5 4.7 5.2 ;
      RECT 2.95 3.5 5.1 3.8 ;
      RECT 4.8 1.55 5.1 3.8 ;
      RECT 2.95 2.75 3.25 3.8 ;
      RECT 2.8 2.75 3.25 3.2 ;
      RECT 4.4 1.55 5.1 1.8 ;
      RECT 4.4 0.95 4.7 1.8 ;
      RECT 2.4 3.5 2.7 5.2 ;
      RECT 2.1 1.55 2.4 3.9 ;
      RECT 2.4 0.95 2.7 1.8 ;
      RECT 1.45 0.95 1.75 5.2 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 5.4 2.85 5.9 3.15 ;
      RECT 4.05 2.8 4.55 3.25 ;
      RECT 3.95 2.05 4.45 2.35 ;
  END
END gf180mcu_osu_sc_gp9t3v3__lshifup
