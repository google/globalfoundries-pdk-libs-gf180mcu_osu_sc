# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__nor2_1 0 0 ;
  SIZE 2.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.8 0.7 ;
        RECT 2.1 0 2.35 1.9 ;
        RECT 0.4 0 0.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 3.6 0.95 3.9 ;
      LAYER Metal2 ;
        RECT 0.45 3.55 0.95 3.95 ;
      LAYER Via1 ;
        RECT 0.57 3.62 0.83 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.85 2.95 2.35 3.25 ;
      LAYER Metal2 ;
        RECT 1.85 2.9 2.35 3.3 ;
      LAYER Via1 ;
        RECT 1.97 2.97 2.23 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 4.85 2.2 7.25 ;
        RECT 1.25 4.85 2.2 5.1 ;
        RECT 1.15 4.25 1.65 4.55 ;
        RECT 1.25 1.05 1.5 5.1 ;
      LAYER Metal2 ;
        RECT 1.15 4.2 1.65 4.6 ;
      LAYER Via1 ;
        RECT 1.27 4.27 1.53 4.53 ;
    END
  END Y
END gf180mcu_osu_sc_gp12t3v3__nor2_1
