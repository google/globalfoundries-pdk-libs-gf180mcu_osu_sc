# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffsrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsrn_1 0 0 ;
  SIZE 20.45 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 20.45 8.3 ;
        RECT 18.8 5.55 19.05 8.3 ;
        RECT 15.5 6.8 15.75 8.3 ;
        RECT 13.9 5.55 14.15 8.3 ;
        RECT 11.3 6.3 11.55 8.3 ;
        RECT 8.5 5.55 8.75 8.3 ;
        RECT 5.45 5.55 5.7 8.3 ;
        RECT 3.85 6.3 4.1 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 20.45 0.7 ;
        RECT 18.8 0 19.05 1.9 ;
        RECT 17.05 0 17.3 1.9 ;
        RECT 14.8 0 15.05 1.9 ;
        RECT 13.9 0 14.15 1.9 ;
        RECT 11.3 0 11.55 1.9 ;
        RECT 8.5 0 8.75 1.5 ;
        RECT 5.45 0 5.7 1.9 ;
        RECT 4.55 0 4.8 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 13.65 2.95 14.15 3.25 ;
      LAYER Metal2 ;
        RECT 13.65 2.9 14.15 3.3 ;
      LAYER Via1 ;
        RECT 13.77 2.97 14.03 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 3.6 6.45 3.9 ;
      LAYER Metal2 ;
        RECT 5.95 3.55 6.45 3.95 ;
      LAYER Via1 ;
        RECT 6.07 3.62 6.33 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 19.65 4.9 20.15 5.25 ;
        RECT 19.65 4.85 20.1 5.25 ;
        RECT 19.65 1.05 19.9 7.25 ;
      LAYER Metal2 ;
        RECT 19.65 4.9 20.15 5.2 ;
        RECT 19.7 4.85 20.1 5.25 ;
      LAYER Via1 ;
        RECT 19.77 4.92 20.03 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17.95 4.25 19.4 4.55 ;
        RECT 19.05 2.15 19.3 4.55 ;
        RECT 17.95 2.15 19.3 2.4 ;
        RECT 17.95 4.25 18.2 7.25 ;
        RECT 17.95 1.05 18.2 2.4 ;
      LAYER Metal2 ;
        RECT 18.9 4.25 19.4 4.55 ;
        RECT 18.95 4.2 19.35 4.6 ;
      LAYER Via1 ;
        RECT 19.02 4.27 19.28 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15.7 4.25 16.2 4.55 ;
        RECT 3.4 4.25 3.9 4.55 ;
      LAYER Metal2 ;
        RECT 15.7 4.2 16.2 4.6 ;
        RECT 3.5 5.55 16.1 5.85 ;
        RECT 15.8 4.2 16.1 5.85 ;
        RECT 3.4 4.2 3.9 4.6 ;
        RECT 3.5 4.2 3.8 5.85 ;
      LAYER Via1 ;
        RECT 3.52 4.27 3.78 4.53 ;
        RECT 15.82 4.27 16.08 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 18.2 2.9 18.6 3.3 ;
      RECT 17.85 2.95 18.65 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 16.6 2.2 17.2 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 16.6 1 16.9 2.6 ;
      RECT 2.75 1 16.9 1.3 ;
      RECT 14.7 2.2 15.2 2.6 ;
      RECT 14.7 1.65 15.1 2.6 ;
      RECT 9.85 1.6 10.25 2 ;
      RECT 9.8 1.65 15.1 1.95 ;
      RECT 14.75 4.85 15.15 5.25 ;
      RECT 10.8 4.85 11.2 5.25 ;
      RECT 10.75 4.9 15.2 5.2 ;
      RECT 12.95 4.2 13.4 4.6 ;
      RECT 11.75 4.2 12.15 4.6 ;
      RECT 10.1 4.2 10.6 4.6 ;
      RECT 7.3 4.2 7.75 4.6 ;
      RECT 7.3 4.25 13.4 4.55 ;
      RECT 12.1 2.9 12.5 3.3 ;
      RECT 10.15 2.9 10.55 3.3 ;
      RECT 10.1 2.95 12.6 3.25 ;
      RECT 10.85 3.55 11.25 3.95 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 8.15 2.25 8.55 2.65 ;
      RECT 4.4 2.25 4.9 2.65 ;
      RECT 4.4 2.3 8.6 2.6 ;
      RECT 17.1 4.85 17.6 5.25 ;
      RECT 4.4 3.55 4.9 3.95 ;
    LAYER Via1 ;
      RECT 18.27 2.97 18.53 3.23 ;
      RECT 17.22 4.92 17.48 5.18 ;
      RECT 16.82 2.27 17.08 2.53 ;
      RECT 14.82 2.27 15.08 2.53 ;
      RECT 14.82 4.92 15.08 5.18 ;
      RECT 13.02 4.27 13.28 4.53 ;
      RECT 12.17 2.97 12.43 3.23 ;
      RECT 11.82 4.27 12.08 4.53 ;
      RECT 10.92 3.62 11.18 3.88 ;
      RECT 10.87 4.92 11.13 5.18 ;
      RECT 10.22 2.97 10.48 3.23 ;
      RECT 10.22 4.27 10.48 4.53 ;
      RECT 9.92 1.67 10.18 1.93 ;
      RECT 8.22 2.32 8.48 2.58 ;
      RECT 7.42 4.27 7.68 4.53 ;
      RECT 4.52 2.32 4.78 2.58 ;
      RECT 4.52 3.62 4.78 3.88 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 17.2 2.95 17.45 7.25 ;
      RECT 14.8 4.8 15.1 5.3 ;
      RECT 14.8 4.9 17.6 5.2 ;
      RECT 16.2 2.95 18.65 3.25 ;
      RECT 16.2 1.05 16.45 3.25 ;
      RECT 16.35 6.3 16.6 7.25 ;
      RECT 14.65 6.3 14.9 7.25 ;
      RECT 14.65 6.3 16.6 6.55 ;
      RECT 13.05 1.05 13.3 7.25 ;
      RECT 13 1.8 13.3 5.65 ;
      RECT 12.95 4.25 13.4 4.55 ;
      RECT 12.15 4.85 12.4 7.25 ;
      RECT 12.15 4.85 12.7 5.1 ;
      RECT 12.45 3.65 12.7 5.1 ;
      RECT 12.15 2.85 12.45 3.9 ;
      RECT 12.15 1.05 12.4 3.9 ;
      RECT 10.75 4.9 11.25 5.2 ;
      RECT 10.85 3.6 11.15 5.2 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 9.55 4.25 10.6 4.55 ;
      RECT 9.55 2.25 9.85 4.55 ;
      RECT 9.45 2.25 9.95 2.55 ;
      RECT 9.9 6.05 10.15 7.25 ;
      RECT 9 6.05 10.15 6.3 ;
      RECT 9 3.55 9.25 6.3 ;
      RECT 8.95 1.7 9.2 3.8 ;
      RECT 8.95 1.7 10.3 1.95 ;
      RECT 9.9 1.65 10.3 1.95 ;
      RECT 9.9 1.05 10.15 1.95 ;
      RECT 8.1 4.9 8.6 5.2 ;
      RECT 8.2 2.3 8.5 5.2 ;
      RECT 8.1 2.3 8.6 2.6 ;
      RECT 6.65 4.25 7.8 4.55 ;
      RECT 7.4 2.3 7.7 4.55 ;
      RECT 7.3 2.3 7.8 2.6 ;
      RECT 7.1 5.05 7.35 7.25 ;
      RECT 5.45 5.05 7.35 5.3 ;
      RECT 5.45 2.35 5.7 5.3 ;
      RECT 4.4 3.6 5.7 3.9 ;
      RECT 5.45 2.35 6.45 2.6 ;
      RECT 6.05 1.65 6.45 2.6 ;
      RECT 6.05 1.65 7.35 1.9 ;
      RECT 7.1 1.05 7.35 1.9 ;
      RECT 4.7 5.8 4.95 7.25 ;
      RECT 3 5.8 3.25 7.25 ;
      RECT 3 5.8 4.95 6.05 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 4.5 2.25 4.75 2.65 ;
      RECT 3.15 2.3 4.9 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 16.7 2.25 17.2 2.55 ;
      RECT 14.7 2.25 15.2 2.55 ;
      RECT 11.7 4.25 12.2 4.55 ;
      RECT 10.1 2.95 10.6 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsrn_1
