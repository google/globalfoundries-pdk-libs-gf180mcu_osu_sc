# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_tinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_tinv_16 0 0 ;
  SIZE 18.3 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 18.3 6.15 ;
        RECT 17.45 3.5 17.7 6.15 ;
        RECT 15.75 3.5 16 6.15 ;
        RECT 14.05 3.5 14.3 6.15 ;
        RECT 12.35 3.5 12.6 6.15 ;
        RECT 10.65 3.5 10.9 6.15 ;
        RECT 8.95 3.5 9.2 6.15 ;
        RECT 7.25 3.5 7.5 6.15 ;
        RECT 5.55 3.5 5.8 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 1.1 3.5 1.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 18.3 0.6 ;
        RECT 17.45 0 17.7 1.8 ;
        RECT 15.75 0 16 1.8 ;
        RECT 14.05 0 14.3 1.8 ;
        RECT 12.35 0 12.6 1.8 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.95 0 9.2 1.8 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.1 0 1.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 1.45 2.25 2.9 ;
      LAYER MET2 ;
        RECT 1.85 1.5 2.35 1.9 ;
      LAYER VIA12 ;
        RECT 1.97 1.57 2.23 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.6 3.5 17.15 3.8 ;
        RECT 16.6 0.95 16.85 5.2 ;
        RECT 4.7 3 16.85 3.25 ;
        RECT 4.7 2.05 16.85 2.3 ;
        RECT 14.9 0.95 15.15 5.2 ;
        RECT 13.2 0.95 13.45 5.2 ;
        RECT 11.5 0.95 11.75 5.2 ;
        RECT 9.8 0.95 10.05 5.2 ;
        RECT 8.1 0.95 8.35 5.2 ;
        RECT 6.4 0.95 6.65 5.2 ;
        RECT 4.7 0.95 4.95 5.2 ;
      LAYER MET2 ;
        RECT 16.65 3.5 17.15 3.8 ;
        RECT 16.7 3.45 17.1 3.85 ;
      LAYER VIA12 ;
        RECT 16.77 3.52 17.03 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.4 2.8 3.95 3.2 ;
    LAYER VIA12 ;
      RECT 3.57 2.87 3.83 3.13 ;
      RECT 2.52 2.87 2.78 3.13 ;
    LAYER MET1 ;
      RECT 3 3.5 3.25 5.2 ;
      RECT 3.05 2.2 3.3 3.7 ;
      RECT 4.15 2.1 4.4 2.55 ;
      RECT 3 0.95 3.25 2.55 ;
      RECT 3 2.2 4.4 2.45 ;
      RECT 2.5 0.95 2.75 5.2 ;
      RECT 2.5 2.75 2.8 3.25 ;
      RECT 3.55 2.75 3.85 3.25 ;
  END
END gf180mcu_osu_sc_9T_tinv_16
