# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_tielo
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_tielo 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 1.55 1.8 1.85 ;
        RECT 1.4 0.95 1.65 1.9 ;
      LAYER MET2 ;
        RECT 1.3 1.5 1.8 1.9 ;
      LAYER VIA12 ;
        RECT 1.42 1.57 1.68 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 2.9 1.65 5.2 ;
      RECT 1.15 2.9 1.65 3.15 ;
  END
END gf180mcu_osu_sc_9T_tielo
