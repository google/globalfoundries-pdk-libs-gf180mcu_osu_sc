* HSPICE file created from gf180mcu_osu_sc_12T_nand2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_nand2_1 A B Y
X0 VDD B Y VDD pmos_3p3 w=34 l=6
X1 Y A VDD VDD pmos_3p3 w=34 l=6
X2 a_28_16 A Y GND nmos_3p3 w=17 l=6
X3 GND B a_28_16 GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
