magic
tech gf180mcuC
timestamp 1661527894
<< nwell >>
rect -17 97 61 159
<< nmos >>
rect 2 55 8 72
rect 19 55 25 72
rect 36 55 42 72
<< pmos >>
rect 2 106 8 140
rect 19 106 25 140
rect 36 106 42 140
<< ndiff >>
rect -8 70 2 72
rect -8 57 -6 70
rect -1 57 2 70
rect -8 55 2 57
rect 8 70 19 72
rect 8 57 11 70
rect 16 57 19 70
rect 8 55 19 57
rect 25 70 36 72
rect 25 57 28 70
rect 33 57 36 70
rect 25 55 36 57
rect 42 70 52 72
rect 42 57 45 70
rect 50 57 52 70
rect 42 55 52 57
<< pdiff >>
rect -8 138 2 140
rect -8 108 -6 138
rect -1 108 2 138
rect -8 106 2 108
rect 8 138 19 140
rect 8 108 11 138
rect 16 108 19 138
rect 8 106 19 108
rect 25 138 36 140
rect 25 113 28 138
rect 33 113 36 138
rect 25 106 36 113
rect 42 138 52 140
rect 42 108 45 138
rect 50 108 52 138
rect 42 106 52 108
<< ndiffc >>
rect -6 57 -1 70
rect 11 57 16 70
rect 28 57 33 70
rect 45 57 50 70
<< pdiffc >>
rect -6 108 -1 138
rect 11 108 16 138
rect 28 113 33 138
rect 45 108 50 138
<< psubdiff >>
rect -8 46 2 48
rect -8 41 -6 46
rect -1 41 2 46
rect -8 39 2 41
rect 16 46 26 48
rect 16 41 18 46
rect 23 41 26 46
rect 16 39 26 41
rect 40 46 50 48
rect 40 41 42 46
rect 47 41 50 46
rect 40 39 50 41
<< nsubdiff >>
rect -8 154 2 156
rect -8 149 -6 154
rect -1 149 2 154
rect -8 147 2 149
rect 16 154 26 156
rect 16 149 18 154
rect 23 149 26 154
rect 16 147 26 149
rect 40 154 50 156
rect 40 149 42 154
rect 47 149 50 154
rect 40 147 50 149
<< psubdiffcont >>
rect -6 41 -1 46
rect 18 41 23 46
rect 42 41 47 46
<< nsubdiffcont >>
rect -6 149 -1 154
rect 18 149 23 154
rect 42 149 47 154
<< polysilicon >>
rect 2 140 8 145
rect 19 140 25 145
rect 36 140 42 145
rect 2 88 8 106
rect 19 104 25 106
rect 36 104 42 106
rect 19 103 42 104
rect 13 101 42 103
rect 13 95 15 101
rect 21 98 42 101
rect 21 95 25 98
rect 13 93 25 95
rect 2 86 14 88
rect 2 80 6 86
rect 12 80 14 86
rect 2 78 14 80
rect 19 80 25 93
rect 2 72 8 78
rect 19 74 42 80
rect 19 72 25 74
rect 36 72 42 74
rect 2 50 8 55
rect 19 50 25 55
rect 36 50 42 55
<< polycontact >>
rect 15 95 21 101
rect 6 80 12 86
<< metal1 >>
rect -17 154 61 159
rect -17 148 -6 154
rect 0 148 18 154
rect 24 148 42 154
rect 48 148 61 154
rect -17 147 61 148
rect -6 138 -1 140
rect -6 101 -1 108
rect 11 138 16 147
rect 28 138 33 140
rect 28 112 33 113
rect 45 138 50 147
rect 11 106 16 108
rect 26 106 28 112
rect 34 106 36 112
rect 45 106 50 108
rect -6 95 15 101
rect 21 95 23 101
rect -6 70 -1 95
rect 4 80 6 86
rect 12 80 14 86
rect -6 55 -1 57
rect 11 70 16 72
rect 11 48 16 57
rect 28 70 33 106
rect 28 55 33 57
rect 45 70 50 72
rect 45 48 50 57
rect -17 47 61 48
rect -17 41 -6 47
rect 0 41 18 47
rect 24 41 42 47
rect 48 41 61 47
rect -17 36 61 41
<< via1 >>
rect -6 149 -1 154
rect -1 149 0 154
rect -6 148 0 149
rect 18 149 23 154
rect 23 149 24 154
rect 18 148 24 149
rect 42 149 47 154
rect 47 149 48 154
rect 42 148 48 149
rect 28 106 34 112
rect 6 80 12 86
rect -6 46 0 47
rect -6 41 -1 46
rect -1 41 0 46
rect 18 46 24 47
rect 18 41 23 46
rect 23 41 24 46
rect 42 46 48 47
rect 42 41 47 46
rect 47 41 48 46
<< metal2 >>
rect -7 154 1 155
rect 17 154 25 155
rect 41 154 49 155
rect -8 148 -6 154
rect 0 148 2 154
rect 16 148 18 154
rect 24 148 26 154
rect 40 148 42 154
rect 48 148 50 154
rect -7 147 1 148
rect 17 147 25 148
rect 41 147 49 148
rect 26 112 36 113
rect 26 106 28 112
rect 34 106 36 112
rect 26 105 36 106
rect 5 86 13 87
rect 4 80 6 86
rect 12 80 14 86
rect 5 79 13 80
rect -7 47 1 48
rect 17 47 25 48
rect 41 47 49 48
rect -8 41 -6 47
rect 0 41 2 47
rect 16 41 18 47
rect 24 41 26 47
rect 40 41 42 47
rect 48 41 50 47
rect -7 40 1 41
rect 17 40 25 41
rect 41 40 49 41
<< labels >>
rlabel metal2 -3 151 -3 151 1 VDD
rlabel metal2 9 83 9 83 1 A
port 1 n
rlabel metal2 -3 44 -3 44 1 GND
rlabel metal2 31 109 31 109 1 Y
port 2 n
<< end >>
