# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_tinv_1 0 0 ;
  SIZE 2.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.8 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 2.2 2.3 2.5 ;
      LAYER MET2 ;
        RECT 1.8 2.15 2.3 2.55 ;
      LAYER VIA12 ;
        RECT 1.92 2.22 2.18 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 4.8 2.3 5.1 ;
      LAYER MET2 ;
        RECT 1.8 4.75 2.3 5.15 ;
      LAYER VIA12 ;
        RECT 1.92 4.82 2.18 5.08 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 5.45 2.2 7.15 ;
        RECT 1.3 1.55 2.2 1.8 ;
        RECT 1.95 0.95 2.2 1.8 ;
        RECT 1.3 5.45 2.2 5.7 ;
        RECT 1.2 3.5 1.7 3.8 ;
        RECT 1.3 1.55 1.55 5.7 ;
      LAYER MET2 ;
        RECT 1.2 3.45 1.7 3.85 ;
      LAYER VIA12 ;
        RECT 1.32 3.52 1.58 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_12T_tinv_1
