# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__and2_1 0 0 ;
  SIZE 4.1 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 4.1 6.35 ;
        RECT 2.25 3.6 2.7 6.35 ;
        RECT 0.55 3.6 0.8 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.1 0.7 ;
        RECT 2.1 0 2.7 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 0.6 2.3 1.1 2.6 ;
        RECT 0.65 2.25 1.05 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 2.95 2.45 3.25 ;
      LAYER Metal2 ;
        RECT 1.95 2.9 2.45 3.3 ;
      LAYER Via1 ;
        RECT 2.07 2.97 2.33 3.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.3 3.6 3.8 3.9 ;
        RECT 3.3 3.55 3.7 3.95 ;
        RECT 3.3 1.05 3.55 5.3 ;
      LAYER Metal2 ;
        RECT 3.3 3.55 3.8 3.95 ;
      LAYER Via1 ;
        RECT 3.42 3.62 3.68 3.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.55 1.65 5.3 ;
      RECT 2.75 2.2 3.05 2.7 ;
      RECT 1.4 2.3 3.05 2.6 ;
      RECT 0.7 1.55 1.65 1.8 ;
      RECT 0.7 1.05 0.95 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__and2_1
