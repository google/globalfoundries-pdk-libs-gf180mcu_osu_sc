
.inc "../../char/techfiles/design.hspice"
.lib "../../char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL GND

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_oai21_1 Y A0 A1 B
X0 Y B a_8_16 GND nmos_3p3 w=17 l=6
X1 GND A0 a_8_16 GND nmos_3p3 w=17 l=6
X2 a_27_106 A0 VDD VDD pmos_3p3 w=34 l=6
X3 VDD B Y VDD pmos_3p3 w=34 l=6
X4 Y A1 a_27_106 VDD pmos_3p3 w=34 l=6
X5 a_8_16 A1 GND GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
