# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xor2_1 0 0 ;
  SIZE 6.7 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 6.7 6.35 ;
        RECT 5 3.9 5.25 6.35 ;
        RECT 1.4 3.9 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 6.7 0.7 ;
        RECT 5 0 5.25 1.85 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.1 2.3 1.6 2.6 ;
      LAYER Metal2 ;
        RECT 1.1 2.3 1.6 2.6 ;
        RECT 1.15 2.25 1.55 2.65 ;
      LAYER Via1 ;
        RECT 1.22 2.32 1.48 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.1 2.3 5.6 2.6 ;
        RECT 2.35 2.1 5.45 2.4 ;
      LAYER Metal2 ;
        RECT 5.1 2.3 5.6 2.6 ;
        RECT 5.15 2.25 5.55 2.65 ;
      LAYER Via1 ;
        RECT 5.22 2.32 5.48 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.05 1.5 3.55 1.8 ;
        RECT 3.15 1.4 3.45 1.85 ;
        RECT 3.2 1.05 3.45 1.85 ;
        RECT 3.05 4.25 3.55 4.55 ;
        RECT 3.2 4.25 3.45 5.3 ;
        RECT 3.15 4.25 3.45 4.65 ;
      LAYER Metal2 ;
        RECT 3.05 1.45 3.55 1.85 ;
        RECT 3.1 4.2 3.5 4.6 ;
        RECT 3.15 1.45 3.45 4.65 ;
      LAYER Via1 ;
        RECT 3.17 4.27 3.43 4.53 ;
        RECT 3.17 1.52 3.43 1.78 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 5.85 1.05 6.1 5.3 ;
      RECT 2.7 3.75 4.7 4 ;
      RECT 4.45 2.65 4.7 4 ;
      RECT 2.7 3.15 3 4 ;
      RECT 4.45 3.2 6.1 3.5 ;
      RECT 2.6 3.15 3.1 3.4 ;
      RECT 4.45 2.65 4.75 3.5 ;
      RECT 4.35 2.65 4.85 2.95 ;
      RECT 0.55 1.05 0.8 5.3 ;
      RECT 3.65 2.65 3.95 3.5 ;
      RECT 0.55 3.1 2.35 3.35 ;
      RECT 2.05 2.65 2.35 3.35 ;
      RECT 2.05 2.65 3.95 2.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xor2_1
