# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_8 0 0 ;
  SIZE 9.05 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 9.05 6.35 ;
        RECT 8.2 3.6 8.45 6.35 ;
        RECT 6.5 3.6 6.75 6.35 ;
        RECT 4.8 3.6 5.05 6.35 ;
        RECT 3.1 3.6 3.35 6.35 ;
        RECT 1.4 3.6 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 9.05 0.7 ;
        RECT 8.2 0 8.45 1.9 ;
        RECT 6.5 0 6.75 1.9 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 3.1 0 3.35 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 2.3 1.55 2.6 ;
      LAYER Metal2 ;
        RECT 1.05 2.3 1.55 2.6 ;
        RECT 1.1 2.25 1.5 2.65 ;
      LAYER Via1 ;
        RECT 1.17 2.32 1.43 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.25 3.6 7.75 3.9 ;
        RECT 7.35 1.05 7.6 5.3 ;
        RECT 2.25 3.05 7.6 3.35 ;
        RECT 2.25 2.15 7.6 2.45 ;
        RECT 5.65 1.05 5.9 5.3 ;
        RECT 3.95 1.05 4.2 5.3 ;
        RECT 2.25 1.05 2.5 5.3 ;
      LAYER Metal2 ;
        RECT 7.25 3.55 7.75 3.95 ;
      LAYER Via1 ;
        RECT 7.37 3.62 7.63 3.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 5.3 ;
      RECT 0.55 3.05 2 3.35 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_8
