magic
tech gf180mcuC
timestamp 1661527508
<< nwell >>
rect 0 100 172 162
<< nmos >>
rect 19 58 25 75
rect 36 58 42 75
rect 53 58 59 75
rect 85 58 91 75
rect 102 58 108 75
rect 124 58 130 75
rect 141 58 147 75
<< pmos >>
rect 19 109 25 143
rect 36 109 42 143
rect 53 109 59 143
rect 85 109 91 143
rect 102 109 108 143
rect 124 109 130 143
rect 141 109 147 143
<< ndiff >>
rect 9 69 19 75
rect 9 60 11 69
rect 16 60 19 69
rect 9 58 19 60
rect 25 73 36 75
rect 25 60 28 73
rect 33 60 36 73
rect 25 58 36 60
rect 42 58 53 75
rect 59 73 69 75
rect 59 60 62 73
rect 67 60 69 73
rect 59 58 69 60
rect 75 66 85 75
rect 75 60 77 66
rect 82 60 85 66
rect 75 58 85 60
rect 91 73 102 75
rect 91 68 94 73
rect 99 68 102 73
rect 91 58 102 68
rect 108 66 124 75
rect 108 60 111 66
rect 116 60 124 66
rect 108 58 124 60
rect 130 73 141 75
rect 130 60 133 73
rect 138 60 141 73
rect 130 58 141 60
rect 147 73 162 75
rect 147 60 155 73
rect 160 60 162 73
rect 147 58 162 60
<< pdiff >>
rect 9 141 19 143
rect 9 116 11 141
rect 16 116 19 141
rect 9 109 19 116
rect 25 141 36 143
rect 25 111 28 141
rect 33 111 36 141
rect 25 109 36 111
rect 42 141 53 143
rect 42 111 45 141
rect 50 111 53 141
rect 42 109 53 111
rect 59 141 69 143
rect 59 111 62 141
rect 67 111 69 141
rect 59 109 69 111
rect 75 141 85 143
rect 75 111 77 141
rect 82 111 85 141
rect 75 109 85 111
rect 91 109 102 143
rect 108 141 124 143
rect 108 111 111 141
rect 121 111 124 141
rect 108 109 124 111
rect 130 141 141 143
rect 130 131 133 141
rect 138 131 141 141
rect 130 109 141 131
rect 147 141 162 143
rect 147 111 150 141
rect 160 111 162 141
rect 147 109 162 111
<< ndiffc >>
rect 11 60 16 69
rect 28 60 33 73
rect 62 60 67 73
rect 77 60 82 66
rect 94 68 99 73
rect 111 60 116 66
rect 133 60 138 73
rect 155 60 160 73
<< pdiffc >>
rect 11 116 16 141
rect 28 111 33 141
rect 45 111 50 141
rect 62 111 67 141
rect 77 111 82 141
rect 111 111 121 141
rect 133 131 138 141
rect 150 111 160 141
<< psubdiff >>
rect 9 49 18 51
rect 9 44 11 49
rect 16 44 18 49
rect 9 42 18 44
rect 33 49 42 51
rect 33 44 35 49
rect 40 44 42 49
rect 33 42 42 44
rect 57 49 66 51
rect 57 44 59 49
rect 64 44 66 49
rect 57 42 66 44
rect 81 49 90 51
rect 81 44 83 49
rect 88 44 90 49
rect 81 42 90 44
rect 105 49 114 51
rect 105 44 107 49
rect 112 44 114 49
rect 105 42 114 44
rect 134 49 143 51
rect 134 44 136 49
rect 141 44 143 49
rect 134 42 143 44
<< nsubdiff >>
rect 9 157 18 159
rect 9 152 11 157
rect 16 152 18 157
rect 9 150 18 152
rect 33 157 42 159
rect 33 152 35 157
rect 40 152 42 157
rect 33 150 42 152
rect 57 157 66 159
rect 57 152 59 157
rect 64 152 66 157
rect 57 150 66 152
rect 81 157 90 159
rect 81 152 83 157
rect 88 152 90 157
rect 81 150 90 152
rect 105 157 114 159
rect 105 152 107 157
rect 112 152 114 157
rect 105 150 114 152
rect 129 157 138 159
rect 129 152 131 157
rect 136 152 138 157
rect 129 150 138 152
<< psubdiffcont >>
rect 11 44 16 49
rect 35 44 40 49
rect 59 44 64 49
rect 83 44 88 49
rect 107 44 112 49
rect 136 44 141 49
<< nsubdiffcont >>
rect 11 152 16 157
rect 35 152 40 157
rect 59 152 64 157
rect 83 152 88 157
rect 107 152 112 157
rect 131 152 136 157
<< polysilicon >>
rect 19 143 25 148
rect 36 143 42 148
rect 53 143 59 148
rect 85 143 91 148
rect 102 143 108 148
rect 124 143 130 148
rect 141 143 147 148
rect 19 106 25 109
rect 19 104 31 106
rect 19 98 23 104
rect 29 98 31 104
rect 19 96 31 98
rect 19 75 25 96
rect 36 91 42 109
rect 30 89 42 91
rect 53 90 59 109
rect 85 91 91 109
rect 30 83 32 89
rect 38 83 42 89
rect 30 81 42 83
rect 36 75 42 81
rect 47 88 59 90
rect 47 82 49 88
rect 55 82 59 88
rect 47 80 59 82
rect 78 89 91 91
rect 78 83 80 89
rect 86 83 91 89
rect 78 81 91 83
rect 53 75 59 80
rect 85 75 91 81
rect 102 87 108 109
rect 124 107 130 109
rect 124 105 136 107
rect 124 99 128 105
rect 134 99 136 105
rect 124 97 136 99
rect 102 85 112 87
rect 102 79 104 85
rect 110 79 112 85
rect 102 77 112 79
rect 102 75 108 77
rect 124 75 130 97
rect 141 91 147 109
rect 135 89 147 91
rect 135 83 137 89
rect 143 83 147 89
rect 135 81 147 83
rect 141 75 147 81
rect 19 53 25 58
rect 36 53 42 58
rect 53 53 59 58
rect 85 53 91 58
rect 102 53 108 58
rect 124 53 130 58
rect 141 53 147 58
<< polycontact >>
rect 23 98 29 104
rect 32 83 38 89
rect 49 82 55 88
rect 80 83 86 89
rect 128 99 134 105
rect 104 79 110 85
rect 137 83 143 89
<< metal1 >>
rect 0 157 172 162
rect 0 151 11 157
rect 17 151 35 157
rect 41 151 59 157
rect 65 151 83 157
rect 89 151 107 157
rect 113 151 131 157
rect 137 151 172 157
rect 0 150 172 151
rect 11 141 16 143
rect 11 115 16 116
rect 28 141 33 150
rect 8 109 10 115
rect 16 109 18 115
rect 28 109 33 111
rect 45 141 50 143
rect 11 69 16 109
rect 45 104 50 111
rect 62 141 67 150
rect 62 109 67 111
rect 77 141 82 150
rect 77 109 82 111
rect 111 141 121 143
rect 133 141 138 150
rect 133 129 138 131
rect 150 141 160 143
rect 111 109 121 111
rect 150 109 160 111
rect 21 98 23 104
rect 29 98 62 104
rect 68 98 70 104
rect 111 99 116 109
rect 126 99 128 105
rect 134 99 136 105
rect 155 103 160 109
rect 155 102 162 103
rect 30 83 32 89
rect 38 83 40 89
rect 47 82 49 88
rect 55 82 57 88
rect 49 76 55 82
rect 11 58 16 60
rect 28 73 33 75
rect 47 70 49 76
rect 55 70 57 76
rect 62 73 67 98
rect 94 94 121 99
rect 154 96 156 102
rect 162 96 164 102
rect 155 95 162 96
rect 78 83 80 89
rect 86 83 88 89
rect 28 51 33 60
rect 94 73 99 94
rect 115 89 135 94
rect 104 85 110 87
rect 130 83 137 89
rect 143 83 145 89
rect 104 77 110 79
rect 133 73 138 75
rect 62 58 67 60
rect 77 66 82 68
rect 94 66 99 68
rect 111 66 116 68
rect 82 60 111 61
rect 77 56 116 60
rect 133 51 138 60
rect 155 73 160 95
rect 155 58 160 60
rect 0 50 172 51
rect 0 44 11 50
rect 17 44 35 50
rect 41 44 59 50
rect 65 44 83 50
rect 89 44 107 50
rect 113 44 136 50
rect 142 44 172 50
rect 0 39 172 44
<< via1 >>
rect 11 152 16 157
rect 16 152 17 157
rect 11 151 17 152
rect 35 152 40 157
rect 40 152 41 157
rect 35 151 41 152
rect 59 152 64 157
rect 64 152 65 157
rect 59 151 65 152
rect 83 152 88 157
rect 88 152 89 157
rect 83 151 89 152
rect 107 152 112 157
rect 112 152 113 157
rect 107 151 113 152
rect 131 152 136 157
rect 136 152 137 157
rect 131 151 137 152
rect 10 109 16 115
rect 62 98 68 104
rect 128 99 134 105
rect 32 83 38 89
rect 49 70 55 76
rect 156 96 162 102
rect 80 83 86 89
rect 104 79 110 85
rect 11 49 17 50
rect 11 44 16 49
rect 16 44 17 49
rect 35 49 41 50
rect 35 44 40 49
rect 40 44 41 49
rect 59 49 65 50
rect 59 44 64 49
rect 64 44 65 49
rect 83 49 89 50
rect 83 44 88 49
rect 88 44 89 49
rect 107 49 113 50
rect 107 44 112 49
rect 112 44 113 49
rect 136 49 142 50
rect 136 44 141 49
rect 141 44 142 49
<< metal2 >>
rect 10 157 18 158
rect 34 157 42 158
rect 58 157 66 158
rect 82 157 90 158
rect 106 157 114 158
rect 130 157 138 158
rect 9 151 11 157
rect 17 151 19 157
rect 33 151 35 157
rect 41 151 43 157
rect 57 151 59 157
rect 65 151 67 157
rect 81 151 83 157
rect 89 151 91 157
rect 105 151 107 157
rect 113 151 115 157
rect 129 151 131 157
rect 137 151 139 157
rect 10 150 18 151
rect 34 150 42 151
rect 58 150 66 151
rect 82 150 90 151
rect 106 150 114 151
rect 130 150 138 151
rect 8 115 18 116
rect 8 109 10 115
rect 16 109 18 115
rect 8 108 18 109
rect 126 105 136 106
rect 60 104 70 105
rect 126 104 128 105
rect 60 98 62 104
rect 68 99 128 104
rect 134 99 136 105
rect 68 98 136 99
rect 154 102 164 103
rect 60 97 70 98
rect 154 96 156 102
rect 162 96 164 102
rect 154 95 164 96
rect 30 89 40 90
rect 78 89 88 90
rect 30 83 32 89
rect 38 83 80 89
rect 86 83 88 89
rect 104 86 110 87
rect 30 82 40 83
rect 78 82 88 83
rect 103 85 111 86
rect 103 79 104 85
rect 110 79 111 85
rect 103 78 111 79
rect 48 76 56 77
rect 103 76 110 78
rect 47 70 49 76
rect 55 70 110 76
rect 48 69 56 70
rect 10 50 18 51
rect 34 50 42 51
rect 58 50 66 51
rect 82 50 90 51
rect 106 50 114 51
rect 135 50 143 51
rect 9 44 11 50
rect 17 44 19 50
rect 33 44 35 50
rect 41 44 43 50
rect 57 44 59 50
rect 65 44 67 50
rect 81 44 83 50
rect 89 44 91 50
rect 105 44 107 50
rect 113 44 115 50
rect 134 44 136 50
rect 142 44 144 50
rect 10 43 18 44
rect 34 43 42 44
rect 58 43 66 44
rect 82 43 90 44
rect 106 43 114 44
rect 135 43 143 44
<< labels >>
rlabel metal2 14 154 14 154 1 VDD
rlabel metal2 35 86 35 86 1 A
port 1 n
rlabel metal2 14 47 14 47 1 GND
rlabel metal2 159 99 159 99 1 S
port 3 n
rlabel metal2 52 73 52 73 1 B
port 5 n
rlabel metal2 12 112 12 112 1 CO
port 4 n
<< end >>
