# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi21_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 1.4 6.2 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.95 0 3.2 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 4.15 2.1 4.45 ;
      LAYER MET2 ;
        RECT 1.6 4.1 2.1 4.5 ;
      LAYER VIA12 ;
        RECT 1.72 4.17 1.98 4.43 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 3.5 2.85 3.8 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.8 3.5 5.1 ;
        RECT 3.1 2.55 3.35 7.15 ;
        RECT 2.1 2.55 3.35 2.8 ;
        RECT 2.1 0.95 2.35 2.8 ;
      LAYER MET2 ;
        RECT 3 4.75 3.5 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 4.82 3.38 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.25 5.7 2.5 7.15 ;
      RECT 0.55 5.7 0.8 7.15 ;
      RECT 0.55 5.7 2.5 5.95 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi21_1
