

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_buf_2 A Y
X0 VDD a_n8_16 Y VDD pmos_3p3 w=34 l=6
X1 Y a_n8_16 VDD VDD pmos_3p3 w=34 l=6
X2 Y a_n8_16 GND GND nmos_3p3 w=17 l=6
X3 VDD A a_n8_16 VDD pmos_3p3 w=34 l=6
X4 GND a_n8_16 Y GND nmos_3p3 w=17 l=6
X5 GND A a_n8_16 GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
