* HSPICE file created from gf180mcu_osu_sc_12T_addh_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/OSU_180/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/OSU_180/char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL GND

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_addh_1 A B S CO
X0 VDD B a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 A VDD VDD pmos_3p3 w=34 l=6
X2 VDD a_19_14 CO VDD pmos_3p3 w=34 l=6
X3 a_19_14 B a_42_19 GND nmos_3p3 w=17 l=6
X4 S a_91_19 GND GND nmos_3p3 w=17 l=6
X5 GND a_19_14 CO GND nmos_3p3 w=17 l=6
X6 S a_91_19 VDD VDD pmos_3p3 w=34 l=6
X7 a_91_19 B a_91_109 VDD pmos_3p3 w=34 l=6
X8 VDD a_19_14 a_91_19 VDD pmos_3p3 w=34 l=6
X9 a_91_109 A VDD VDD pmos_3p3 w=34 l=6
X10 a_91_19 A a_75_19 GND nmos_3p3 w=17 l=6
X11 a_42_19 A GND GND nmos_3p3 w=17 l=6
X12 GND a_19_14 a_75_19 GND nmos_3p3 w=17 l=6
X13 a_75_19 B a_91_19 GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
