magic
tech gf180mcuC
timestamp 1661875506
<< nwell >>
rect 0 61 128 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 49 19 55 36
rect 72 19 78 36
rect 85 19 91 36
rect 102 19 108 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 49 70 55 104
rect 72 70 78 104
rect 85 70 91 104
rect 102 70 108 104
<< ndiff >>
rect 58 36 68 37
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 19 49 36
rect 55 35 72 36
rect 55 21 61 35
rect 66 21 72 35
rect 55 19 72 21
rect 78 19 85 36
rect 91 34 102 36
rect 91 21 94 34
rect 99 21 102 34
rect 91 19 102 21
rect 108 34 118 36
rect 108 21 111 34
rect 116 21 118 34
rect 108 19 118 21
<< pdiff >>
rect 9 102 19 104
rect 9 94 11 102
rect 16 94 19 102
rect 9 70 19 94
rect 25 102 36 104
rect 25 94 28 102
rect 33 94 36 102
rect 25 70 36 94
rect 42 70 49 104
rect 55 102 72 104
rect 55 94 61 102
rect 66 94 72 102
rect 55 70 72 94
rect 78 70 85 104
rect 91 102 102 104
rect 91 94 94 102
rect 99 94 102 102
rect 91 70 102 94
rect 108 102 118 104
rect 108 94 111 102
rect 116 94 118 102
rect 108 70 118 94
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 61 21 66 35
rect 94 21 99 34
rect 111 21 116 34
<< pdiffc >>
rect 11 94 16 102
rect 28 94 33 102
rect 61 94 66 102
rect 94 94 99 102
rect 111 94 116 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
rect 81 118 90 120
rect 81 113 83 118
rect 88 113 90 118
rect 81 111 90 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
rect 107 113 112 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 49 104 55 109
rect 72 104 78 109
rect 85 104 91 109
rect 102 104 108 109
rect 19 52 25 70
rect 36 68 42 70
rect 31 66 42 68
rect 31 60 33 66
rect 39 60 42 66
rect 31 58 42 60
rect 49 68 55 70
rect 72 68 78 70
rect 85 68 91 70
rect 102 68 108 70
rect 49 66 63 68
rect 49 60 55 66
rect 61 60 63 66
rect 49 58 63 60
rect 70 66 80 68
rect 70 60 72 66
rect 78 60 80 66
rect 85 63 108 68
rect 70 58 80 60
rect 19 50 35 52
rect 19 44 27 50
rect 33 49 35 50
rect 33 44 42 49
rect 19 42 42 44
rect 19 36 25 42
rect 36 36 42 42
rect 49 36 55 58
rect 102 52 108 63
rect 60 50 70 52
rect 91 50 108 52
rect 60 44 62 50
rect 68 44 78 50
rect 91 47 93 50
rect 60 42 78 44
rect 72 36 78 42
rect 85 44 93 47
rect 99 44 108 50
rect 85 42 108 44
rect 85 36 91 42
rect 102 36 108 42
rect 19 14 25 19
rect 36 14 42 19
rect 49 14 55 19
rect 72 14 78 19
rect 85 14 91 19
rect 102 14 108 19
<< polycontact >>
rect 33 60 39 66
rect 55 60 61 66
rect 72 60 78 66
rect 27 44 33 50
rect 62 44 68 50
rect 93 44 99 50
<< metal1 >>
rect 0 118 128 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 128 118
rect 0 111 128 112
rect 11 102 16 104
rect 11 66 16 94
rect 28 102 33 111
rect 61 102 66 104
rect 28 92 33 94
rect 60 94 61 95
rect 60 89 66 94
rect 94 102 99 111
rect 94 92 99 94
rect 111 102 116 104
rect 60 81 66 83
rect 111 76 116 94
rect 55 71 116 76
rect 55 66 61 71
rect 11 60 33 66
rect 39 60 48 66
rect 11 34 16 60
rect 42 50 48 60
rect 70 60 72 66
rect 78 60 80 66
rect 55 58 61 60
rect 25 44 27 50
rect 33 44 35 50
rect 42 44 62 50
rect 68 44 70 50
rect 91 44 93 50
rect 99 44 101 50
rect 60 37 66 39
rect 11 19 16 21
rect 28 34 33 36
rect 60 28 61 31
rect 28 12 33 21
rect 61 19 66 21
rect 94 34 99 36
rect 94 12 99 21
rect 111 34 116 71
rect 111 19 116 21
rect 0 11 128 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 128 11
rect 0 0 128 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 60 83 66 89
rect 72 60 78 66
rect 27 44 33 50
rect 93 44 99 50
rect 60 35 66 37
rect 60 31 61 35
rect 61 31 66 35
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 60 90 66 95
rect 59 89 67 90
rect 59 83 60 89
rect 66 83 67 89
rect 59 82 67 83
rect 59 81 66 82
rect 27 51 33 52
rect 26 50 34 51
rect 26 44 27 50
rect 33 44 34 50
rect 26 43 34 44
rect 27 24 33 43
rect 59 38 65 81
rect 72 67 79 68
rect 71 66 80 67
rect 71 60 72 66
rect 78 60 80 66
rect 71 59 80 60
rect 72 58 80 59
rect 58 37 68 38
rect 58 31 60 37
rect 66 31 68 37
rect 58 30 68 31
rect 74 24 80 58
rect 93 51 99 52
rect 92 50 100 51
rect 91 44 93 50
rect 99 44 101 50
rect 92 43 100 44
rect 93 42 99 43
rect 27 18 80 24
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 30 47 30 47 1 A
port 1 n
rlabel metal2 96 47 96 47 1 B
port 4 n
rlabel metal2 63 85 63 85 1 Y
port 3 n
<< end >>
