# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_clkinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_clkinv_8 0 0 ;
  SIZE 8.15 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 8.15 8.1 ;
        RECT 7.35 5.45 7.6 8.1 ;
        RECT 5.65 5.45 5.9 8.1 ;
        RECT 3.95 5.45 4.2 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
      LAYER MET2 ;
        RECT 6.45 7.55 6.95 7.85 ;
        RECT 6.5 7.5 6.9 7.9 ;
        RECT 5.25 7.55 5.75 7.85 ;
        RECT 5.3 7.5 5.7 7.9 ;
        RECT 4.05 7.55 4.55 7.85 ;
        RECT 4.1 7.5 4.5 7.9 ;
        RECT 2.85 7.55 3.35 7.85 ;
        RECT 2.9 7.5 3.3 7.9 ;
        RECT 1.65 7.55 2.15 7.85 ;
        RECT 1.7 7.5 2.1 7.9 ;
        RECT 0.45 7.55 0.95 7.85 ;
        RECT 0.5 7.5 0.9 7.9 ;
      LAYER VIA12 ;
        RECT 0.57 7.57 0.83 7.83 ;
        RECT 1.77 7.57 2.03 7.83 ;
        RECT 2.97 7.57 3.23 7.83 ;
        RECT 4.17 7.57 4.43 7.83 ;
        RECT 5.37 7.57 5.63 7.83 ;
        RECT 6.57 7.57 6.83 7.83 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.15 0.6 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
      LAYER MET2 ;
        RECT 6.45 0.25 6.95 0.55 ;
        RECT 6.5 0.2 6.9 0.6 ;
        RECT 5.25 0.25 5.75 0.55 ;
        RECT 5.3 0.2 5.7 0.6 ;
        RECT 4.05 0.25 4.55 0.55 ;
        RECT 4.1 0.2 4.5 0.6 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
        RECT 4.17 0.27 4.43 0.53 ;
        RECT 5.37 0.27 5.63 0.53 ;
        RECT 6.57 0.27 6.83 0.53 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.5 0.95 6.75 7.15 ;
        RECT 1.4 4.45 6.75 4.7 ;
        RECT 6.35 4.35 6.75 4.7 ;
        RECT 1.4 2.05 6.75 2.3 ;
        RECT 4.8 0.95 5.05 7.15 ;
        RECT 3.1 0.95 3.35 7.15 ;
        RECT 1.4 0.95 1.65 7.15 ;
      LAYER MET2 ;
        RECT 6.35 4.35 6.85 4.75 ;
      LAYER VIA12 ;
        RECT 6.47 4.42 6.73 4.68 ;
    END
  END Y
END gf180mcu_osu_sc_12T_clkinv_8
