magic
tech gf180mcuC
timestamp 1660768231
<< nwell >>
rect 0 97 56 159
<< nmos >>
rect 16 55 22 72
rect 33 55 39 72
<< pmos >>
rect 19 106 25 140
rect 30 106 36 140
<< ndiff >>
rect 6 70 16 72
rect 6 57 8 70
rect 13 57 16 70
rect 6 55 16 57
rect 22 70 33 72
rect 22 57 25 70
rect 30 57 33 70
rect 22 55 33 57
rect 39 70 49 72
rect 39 57 42 70
rect 47 57 49 70
rect 39 55 49 57
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 106 30 140
rect 36 138 46 140
rect 36 115 39 138
rect 44 115 46 138
rect 36 106 46 115
<< ndiffc >>
rect 8 57 13 70
rect 25 57 30 70
rect 42 57 47 70
<< pdiffc >>
rect 11 108 16 138
rect 39 115 44 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
<< polysilicon >>
rect 19 140 25 145
rect 30 140 36 145
rect 19 102 25 106
rect 16 97 25 102
rect 30 103 36 106
rect 30 101 39 103
rect 30 99 47 101
rect 30 97 39 99
rect 16 88 22 97
rect 8 86 22 88
rect 8 80 11 86
rect 17 80 22 86
rect 8 78 22 80
rect 16 72 22 78
rect 33 93 39 97
rect 45 93 47 99
rect 33 91 47 93
rect 33 72 39 91
rect 16 50 22 55
rect 33 50 39 55
<< polycontact >>
rect 11 80 17 86
rect 39 93 45 99
<< metal1 >>
rect 0 154 56 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 56 154
rect 0 147 56 148
rect 11 138 16 147
rect 39 138 44 140
rect 39 113 44 115
rect 25 112 44 113
rect 11 106 16 108
rect 23 106 25 112
rect 31 108 44 112
rect 31 106 33 108
rect 9 80 11 86
rect 17 80 19 86
rect 8 70 13 72
rect 8 48 13 57
rect 25 70 30 106
rect 37 93 39 99
rect 45 93 47 99
rect 25 55 30 57
rect 42 70 47 72
rect 42 48 47 57
rect 0 47 56 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 56 47
rect 0 36 56 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 25 106 31 112
rect 11 80 17 86
rect 39 93 45 99
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 10 147 18 148
rect 34 147 42 148
rect 23 112 33 113
rect 23 106 25 112
rect 31 106 33 112
rect 23 105 33 106
rect 37 99 47 100
rect 37 93 39 99
rect 45 93 47 99
rect 37 92 47 93
rect 9 86 19 87
rect 9 80 11 86
rect 17 80 19 86
rect 9 79 19 80
rect 10 47 18 48
rect 34 47 42 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 10 40 18 41
rect 34 40 42 41
<< labels >>
rlabel metal2 13 151 13 151 1 VDD
rlabel metal2 14 44 14 44 1 GND
rlabel metal2 14 83 14 83 1 A
port 1 n
rlabel metal2 28 109 28 109 1 Y
port 2 n
rlabel metal2 42 96 42 96 1 B
port 3 n
<< end >>
