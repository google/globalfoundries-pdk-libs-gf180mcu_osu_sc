VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_tiehi
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_tiehi 0 -0.15 ;
  SIZE 2.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 2.2 7.95 ;
        RECT 0.55 5.3 0.8 7.95 ;
      LAYER MET2 ;
        RECT 0.45 7.4 0.95 7.7 ;
        RECT 0.5 7.35 0.9 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 2.2 0.45 ;
        RECT 0.55 -0.15 0.8 1.65 ;
      LAYER MET2 ;
        RECT 0.45 0.1 0.95 0.4 ;
        RECT 0.5 0.05 0.9 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 4.65 1.8 4.95 ;
        RECT 1.4 4.6 1.65 7 ;
      LAYER MET2 ;
        RECT 1.3 4.6 1.8 5 ;
      LAYER VIA12 ;
        RECT 1.42 4.67 1.68 4.93 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.15 2.05 1.65 2.3 ;
      RECT 1.4 0.8 1.65 2.3 ;
  END
END gf180mcu_osu_sc_12T_tiehi
