# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__lshifdown
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__lshifdown 0 0 ;
  SIZE 4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 2.15 5.55 4 6.15 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 1.85 6.15 ;
        RECT 0.55 3.5 0.85 6.15 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4 0.6 ;
        RECT 2.25 0 2.55 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 0.55 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 2.2 3.5 2.5 ;
        RECT 3.15 0.95 3.45 5.2 ;
      LAYER MET2 ;
        RECT 3.05 2.15 3.55 2.55 ;
      LAYER VIA12 ;
        RECT 3.17 2.22 3.43 2.48 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.3 2.8 2.8 3.2 ;
      RECT 1.45 2.85 2.8 3.15 ;
      RECT 1.45 2.15 1.75 3.15 ;
      RECT 1.35 2.15 1.85 2.55 ;
    LAYER VIA12 ;
      RECT 2.42 2.87 2.68 3.13 ;
      RECT 1.47 2.22 1.73 2.48 ;
    LAYER MET1 ;
      RECT 1.45 0.95 1.75 5.2 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 2.3 2.85 2.8 3.15 ;
      RECT 2.25 3.5 2.55 5.2 ;
  END
END gf180mcu_osu_sc_gp9t3v3__lshifdown
