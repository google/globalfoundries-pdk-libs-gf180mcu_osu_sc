* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffn_1 Q QN D CLK VDD VSS
X0 a_75_109# a_52_14# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# a_52_81# a_42_109# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_131_19# a_52_14# a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X3 a_42_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_75_19# a_52_81# a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X6 VDD a_135_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X7 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X9 VSS a_135_68# a_131_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 a_19_14# a_52_14# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_135_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X13 a_52_14# a_52_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD a_135_68# a_131_109# VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS CLK a_52_81# VSS nmos_3p3 w=0.85u l=0.3u
X16 a_131_109# a_52_81# a_114_19# VDD pmos_3p3 w=1.7u l=0.3u
X17 a_114_19# a_52_14# a_103_109# VDD pmos_3p3 w=1.7u l=0.3u
X18 a_135_68# a_114_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 a_114_19# a_52_81# a_103_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_52_14# a_52_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X21 a_103_109# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD a_9_19# a_75_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_103_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 a_135_68# a_114_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X26 VDD CLK a_52_81# VDD pmos_3p3 w=1.7u l=0.3u
X27 VSS a_9_19# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
