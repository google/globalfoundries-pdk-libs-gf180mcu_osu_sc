VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_or2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_or2_1 0 -0.15 ;
  SIZE 3.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 3.35 1.4 3.65 ;
      LAYER MET2 ;
        RECT 0.9 3.3 1.4 3.7 ;
      LAYER VIA12 ;
        RECT 1.02 3.37 1.28 3.63 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.7 2.15 3 ;
      LAYER MET2 ;
        RECT 1.65 2.65 2.15 3.05 ;
      LAYER VIA12 ;
        RECT 1.77 2.72 2.03 2.98 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 3.8 7.95 ;
        RECT 1.95 5.3 2.35 7.95 ;
      LAYER MET2 ;
        RECT 2.85 7.35 3.35 7.75 ;
        RECT 1.65 7.35 2.15 7.75 ;
        RECT 0.45 7.35 0.95 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
        RECT 1.77 7.42 2.03 7.68 ;
        RECT 2.97 7.42 3.23 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 3.8 0.45 ;
        RECT 2.1 -0.15 2.35 1.65 ;
        RECT 0.4 -0.15 0.65 1.65 ;
      LAYER MET2 ;
        RECT 2.85 0.05 3.35 0.45 ;
        RECT 1.65 0.05 2.15 0.45 ;
        RECT 0.45 0.05 0.95 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
        RECT 1.77 0.12 2.03 0.38 ;
        RECT 2.97 0.12 3.23 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 4.65 3.45 4.95 ;
        RECT 2.95 0.8 3.2 7 ;
      LAYER MET2 ;
        RECT 2.95 4.6 3.45 5 ;
      LAYER VIA12 ;
        RECT 3.07 4.67 3.33 4.93 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.2 3.95 2.7 4.35 ;
    LAYER VIA12 ;
      RECT 2.32 4.02 2.58 4.28 ;
    LAYER MET1 ;
      RECT 0.55 5.1 0.8 7 ;
      RECT 0.4 2.05 0.65 5.35 ;
      RECT 0.4 4 2.7 4.3 ;
      RECT 0.4 2.05 1.5 2.3 ;
      RECT 1.25 0.8 1.5 2.3 ;
  END
END gf180mcu_osu_sc_12T_or2_1
