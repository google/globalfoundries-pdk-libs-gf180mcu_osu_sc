magic
tech gf180mcuC
timestamp 1664894556
<< nwell >>
rect -155 100 25 162
<< nmos >>
rect -135 19 -129 36
rect -115 19 -109 36
rect -101 19 -95 36
rect -84 19 -78 36
rect -70 19 -64 36
rect -50 19 -44 36
rect -18 19 -12 36
rect -1 19 5 36
<< pmos >>
rect -135 109 -129 143
rect -118 109 -112 143
rect -101 109 -95 143
rect -84 109 -78 143
rect -67 109 -61 143
rect -50 109 -44 143
rect -18 109 -12 143
rect -1 109 5 143
<< ndiff >>
rect -145 34 -135 36
rect -145 21 -143 34
rect -138 21 -135 34
rect -145 19 -135 21
rect -129 34 -115 36
rect -129 21 -126 34
rect -118 21 -115 34
rect -129 19 -115 21
rect -109 19 -101 36
rect -95 34 -84 36
rect -95 21 -92 34
rect -87 21 -84 34
rect -95 19 -84 21
rect -78 19 -70 36
rect -64 34 -50 36
rect -64 21 -61 34
rect -53 21 -50 34
rect -64 19 -50 21
rect -44 34 -34 36
rect -44 21 -41 34
rect -36 21 -34 34
rect -44 19 -34 21
rect -28 34 -18 36
rect -28 21 -26 34
rect -21 21 -18 34
rect -28 19 -18 21
rect -12 34 -1 36
rect -12 21 -9 34
rect -4 21 -1 34
rect -12 19 -1 21
rect 5 34 15 36
rect 5 21 8 34
rect 13 21 15 34
rect 5 19 15 21
<< pdiff >>
rect -145 141 -135 143
rect -145 111 -143 141
rect -138 111 -135 141
rect -145 109 -135 111
rect -129 141 -118 143
rect -129 127 -126 141
rect -121 127 -118 141
rect -129 109 -118 127
rect -112 109 -101 143
rect -95 141 -84 143
rect -95 111 -92 141
rect -87 111 -84 141
rect -95 109 -84 111
rect -78 109 -67 143
rect -61 141 -50 143
rect -61 111 -58 141
rect -53 111 -50 141
rect -61 109 -50 111
rect -44 141 -34 143
rect -44 111 -41 141
rect -36 111 -34 141
rect -44 109 -34 111
rect -28 141 -18 143
rect -28 111 -26 141
rect -21 111 -18 141
rect -28 109 -18 111
rect -12 141 -1 143
rect -12 111 -9 141
rect -4 111 -1 141
rect -12 109 -1 111
rect 5 141 15 143
rect 5 111 8 141
rect 13 111 15 141
rect 5 109 15 111
<< ndiffc >>
rect -143 21 -138 34
rect -126 21 -118 34
rect -92 21 -87 34
rect -61 21 -53 34
rect -41 21 -36 34
rect -26 21 -21 34
rect -9 21 -4 34
rect 8 21 13 34
<< pdiffc >>
rect -143 111 -138 141
rect -126 127 -121 141
rect -92 111 -87 141
rect -58 111 -53 141
rect -41 111 -36 141
rect -26 111 -21 141
rect -9 111 -4 141
rect 8 111 13 141
<< psubdiff >>
rect -146 10 -137 12
rect -146 5 -144 10
rect -139 5 -137 10
rect -146 3 -137 5
rect -121 10 -112 12
rect -121 5 -119 10
rect -114 5 -112 10
rect -121 3 -112 5
rect -98 10 -89 12
rect -98 5 -96 10
rect -91 5 -89 10
rect -98 3 -89 5
rect -74 10 -65 12
rect -74 5 -72 10
rect -67 5 -65 10
rect -74 3 -65 5
rect -49 10 -40 12
rect -49 5 -47 10
rect -42 5 -40 10
rect -49 3 -40 5
rect -26 10 -16 12
rect -26 5 -24 10
rect -19 5 -16 10
rect -26 3 -16 5
rect -2 10 7 12
rect -2 5 0 10
rect 5 5 7 10
rect -2 3 7 5
<< nsubdiff >>
rect -146 157 -137 159
rect -146 152 -144 157
rect -139 152 -137 157
rect -146 150 -137 152
rect -121 157 -112 159
rect -121 152 -119 157
rect -114 152 -112 157
rect -121 150 -112 152
rect -98 157 -89 159
rect -98 152 -96 157
rect -91 152 -89 157
rect -98 150 -89 152
rect -74 157 -65 159
rect -74 152 -72 157
rect -67 152 -65 157
rect -74 150 -65 152
rect -49 157 -40 159
rect -49 152 -47 157
rect -42 152 -40 157
rect -49 150 -40 152
rect -25 157 -16 159
rect -25 152 -23 157
rect -18 152 -16 157
rect -25 150 -16 152
rect -1 157 8 159
rect -1 152 1 157
rect 6 152 8 157
rect -1 150 8 152
<< psubdiffcont >>
rect -144 5 -139 10
rect -119 5 -114 10
rect -96 5 -91 10
rect -72 5 -67 10
rect -47 5 -42 10
rect -24 5 -19 10
rect 0 5 5 10
<< nsubdiffcont >>
rect -144 152 -139 157
rect -119 152 -114 157
rect -96 152 -91 157
rect -72 152 -67 157
rect -47 152 -42 157
rect -23 152 -18 157
rect 1 152 6 157
<< polysilicon >>
rect -135 143 -129 148
rect -118 143 -112 148
rect -101 143 -95 148
rect -84 143 -78 148
rect -67 143 -61 148
rect -50 143 -44 148
rect -18 143 -12 148
rect -1 143 5 148
rect -135 91 -129 109
rect -118 91 -112 109
rect -101 102 -95 109
rect -103 100 -93 102
rect -103 94 -101 100
rect -95 94 -93 100
rect -103 92 -93 94
rect -84 91 -78 109
rect -135 89 -123 91
rect -135 83 -132 89
rect -126 83 -123 89
rect -135 81 -123 83
rect -118 89 -108 91
rect -118 83 -116 89
rect -110 83 -108 89
rect -118 81 -108 83
rect -86 89 -76 91
rect -86 83 -84 89
rect -78 83 -76 89
rect -86 81 -76 83
rect -135 36 -129 81
rect -118 45 -112 81
rect -84 70 -78 81
rect -101 64 -78 70
rect -67 78 -61 109
rect -50 91 -44 109
rect -51 89 -41 91
rect -51 83 -49 89
rect -43 83 -41 89
rect -51 81 -41 83
rect -67 76 -55 78
rect -67 70 -63 76
rect -57 70 -55 76
rect -67 68 -55 70
rect -118 41 -109 45
rect -115 36 -109 41
rect -101 36 -95 64
rect -86 57 -76 59
rect -86 51 -84 57
rect -78 51 -76 57
rect -86 49 -76 51
rect -84 36 -78 49
rect -67 45 -61 68
rect -70 41 -61 45
rect -70 36 -64 41
rect -50 36 -44 81
rect -18 78 -12 109
rect -1 91 5 109
rect -7 89 5 91
rect -7 83 -5 89
rect 1 83 5 89
rect -7 81 5 83
rect -20 76 -11 78
rect -20 71 -18 76
rect -13 71 -11 76
rect -20 69 -11 71
rect -18 36 -12 69
rect -1 36 5 81
rect -135 14 -129 19
rect -115 14 -109 19
rect -101 14 -95 19
rect -84 14 -78 19
rect -70 14 -64 19
rect -50 14 -44 19
rect -18 14 -12 19
rect -1 14 5 19
<< polycontact >>
rect -101 94 -95 100
rect -132 83 -126 89
rect -116 83 -110 89
rect -84 83 -78 89
rect -49 83 -43 89
rect -63 70 -57 76
rect -84 51 -78 57
rect -5 83 1 89
rect -18 71 -13 76
<< metal1 >>
rect -155 157 25 162
rect -155 151 -144 157
rect -138 151 -120 157
rect -114 151 -96 157
rect -90 151 -72 157
rect -66 151 -48 157
rect -42 151 -24 157
rect -18 151 0 157
rect 6 151 25 157
rect -155 150 25 151
rect -143 141 -138 143
rect -126 141 -121 150
rect -126 125 -121 127
rect -92 141 -87 143
rect -143 77 -138 111
rect -132 111 -92 114
rect -132 109 -87 111
rect -58 141 -53 150
rect -58 109 -53 111
rect -41 141 -36 143
rect -41 110 -36 111
rect -26 141 -21 143
rect -132 89 -127 109
rect -41 105 -31 110
rect -103 94 -101 100
rect -95 94 -93 100
rect -133 83 -132 89
rect -126 83 -124 89
rect -118 83 -116 89
rect -110 83 -108 89
rect -145 76 -138 77
rect -148 70 -146 76
rect -140 70 -138 76
rect -146 69 -138 70
rect -143 34 -138 69
rect -132 46 -127 83
rect -101 57 -95 94
rect -86 83 -84 89
rect -78 83 -76 89
rect -51 83 -49 89
rect -43 83 -41 89
rect -65 70 -63 76
rect -57 70 -55 76
rect -36 57 -31 105
rect -26 106 -21 111
rect -9 141 -4 150
rect -9 109 -4 111
rect 8 141 13 143
rect -26 102 -18 106
rect 8 103 13 111
rect 8 102 16 103
rect -26 96 -24 102
rect -18 101 -16 102
rect -18 96 1 101
rect -26 95 -18 96
rect -5 89 1 96
rect -20 70 -18 76
rect -12 70 -10 76
rect -101 51 -84 57
rect -78 51 -31 57
rect -132 41 -87 46
rect -36 44 -31 51
rect -5 46 1 83
rect -143 19 -138 21
rect -126 34 -118 36
rect -126 12 -118 21
rect -92 34 -87 41
rect -41 39 -31 44
rect -26 41 1 46
rect 8 96 10 102
rect 16 96 18 102
rect 8 95 16 96
rect -92 19 -87 21
rect -61 34 -53 36
rect -61 12 -53 21
rect -41 34 -36 39
rect -41 19 -36 21
rect -26 34 -21 41
rect -26 19 -21 21
rect -9 34 -4 36
rect -9 12 -4 21
rect 8 34 13 95
rect 8 19 13 21
rect -155 11 25 12
rect -155 5 -144 11
rect -138 5 -120 11
rect -114 5 -96 11
rect -90 5 -72 11
rect -66 5 -48 11
rect -42 5 -24 11
rect -18 5 0 11
rect 6 5 25 11
rect -155 0 25 5
<< via1 >>
rect -144 152 -139 157
rect -139 152 -138 157
rect -144 151 -138 152
rect -120 152 -119 157
rect -119 152 -114 157
rect -120 151 -114 152
rect -96 152 -91 157
rect -91 152 -90 157
rect -96 151 -90 152
rect -72 152 -67 157
rect -67 152 -66 157
rect -72 151 -66 152
rect -48 152 -47 157
rect -47 152 -42 157
rect -48 151 -42 152
rect -24 152 -23 157
rect -23 152 -18 157
rect -24 151 -18 152
rect 0 152 1 157
rect 1 152 6 157
rect 0 151 6 152
rect -116 83 -110 89
rect -146 70 -140 76
rect -84 83 -78 89
rect -49 83 -43 89
rect -63 70 -57 76
rect -24 96 -18 102
rect -18 71 -13 76
rect -13 71 -12 76
rect -18 70 -12 71
rect 10 96 16 102
rect -144 10 -138 11
rect -144 5 -139 10
rect -139 5 -138 10
rect -120 10 -114 11
rect -120 5 -119 10
rect -119 5 -114 10
rect -96 10 -90 11
rect -96 5 -91 10
rect -91 5 -90 10
rect -72 10 -66 11
rect -72 5 -67 10
rect -67 5 -66 10
rect -48 10 -42 11
rect -48 5 -47 10
rect -47 5 -42 10
rect -24 10 -18 11
rect -24 5 -19 10
rect -19 5 -18 10
rect 0 10 6 11
rect 0 5 5 10
rect 5 5 6 10
<< metal2 >>
rect -145 157 -137 158
rect -121 157 -113 158
rect -97 157 -89 158
rect -73 157 -65 158
rect -49 157 -41 158
rect -25 157 -17 158
rect -1 157 7 158
rect -146 151 -144 157
rect -138 151 -136 157
rect -122 151 -120 157
rect -114 151 -112 157
rect -98 151 -96 157
rect -90 151 -88 157
rect -74 151 -72 157
rect -66 151 -64 157
rect -50 151 -48 157
rect -42 151 -40 157
rect -26 151 -24 157
rect -18 151 -16 157
rect -2 151 0 157
rect 6 151 8 157
rect -145 150 -137 151
rect -121 150 -113 151
rect -97 150 -89 151
rect -73 150 -65 151
rect -49 150 -41 151
rect -25 150 -17 151
rect -1 150 7 151
rect -25 102 -17 103
rect 9 102 17 103
rect -26 96 -24 102
rect -18 96 -16 102
rect 8 96 10 102
rect 16 96 18 102
rect -25 95 -17 96
rect 9 95 17 96
rect -118 89 -108 90
rect -85 89 -77 90
rect -51 89 -41 90
rect -118 83 -116 89
rect -110 83 -108 89
rect -86 83 -84 89
rect -78 83 -49 89
rect -43 83 -41 89
rect -118 82 -108 83
rect -85 82 -77 83
rect -51 82 -41 83
rect -148 76 -138 77
rect -64 76 -56 77
rect -20 76 -10 77
rect -148 70 -146 76
rect -140 70 -63 76
rect -57 70 -18 76
rect -12 70 -10 76
rect -148 69 -138 70
rect -64 69 -56 70
rect -20 69 -10 70
rect -145 11 -137 12
rect -121 11 -113 12
rect -97 11 -89 12
rect -73 11 -65 12
rect -49 11 -41 12
rect -25 11 -17 12
rect -1 11 7 12
rect -146 5 -144 11
rect -138 5 -136 11
rect -122 5 -120 11
rect -114 5 -112 11
rect -98 5 -96 11
rect -90 5 -88 11
rect -74 5 -72 11
rect -66 5 -64 11
rect -50 5 -48 11
rect -42 5 -40 11
rect -26 5 -24 11
rect -18 5 -16 11
rect -2 5 0 11
rect 6 5 8 11
rect -145 4 -137 5
rect -121 4 -113 5
rect -97 4 -89 5
rect -73 4 -65 5
rect -49 4 -41 5
rect -25 4 -17 5
rect -1 4 7 5
<< labels >>
rlabel metal2 -141 154 -141 154 1 VDD
rlabel metal2 -141 8 -141 8 1 GND
rlabel metal2 -113 86 -113 86 1 D
port 1 n
rlabel metal2 13 99 13 99 1 Q
port 4 n
rlabel metal2 -81 86 -81 86 1 CLKN
port 5 n
<< end >>
