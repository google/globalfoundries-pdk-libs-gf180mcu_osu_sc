# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__lshifup 0 0 ;
  SIZE 8.15 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.3 6.15 ;
        RECT 0.55 3.5 0.85 6.15 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.9 5.55 8.15 6.15 ;
        RECT 6.4 3.5 6.7 6.15 ;
        RECT 4.35 4.05 4.85 6.15 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.15 0.6 ;
        RECT 6.4 0 6.7 1.8 ;
        RECT 4.35 0 4.85 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.7 2.05 4.2 2.35 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 3.7 2.05 4.2 2.35 ;
        RECT 3.7 2 4.15 2.4 ;
        RECT 3.85 1.4 4.15 2.4 ;
        RECT 0.7 1.4 4.15 1.7 ;
        RECT 0.55 2.15 1.05 2.55 ;
        RECT 0.7 1.4 1 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
        RECT 3.82 2.07 4.08 2.33 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 2.2 7.65 2.5 ;
        RECT 7.3 0.95 7.6 5.2 ;
      LAYER MET2 ;
        RECT 7.2 2.15 7.7 2.55 ;
      LAYER VIA12 ;
        RECT 7.32 2.22 7.58 2.48 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 3.25 3.5 3.75 3.9 ;
      RECT 3.25 3.5 5.5 3.85 ;
      RECT 5.2 2.8 5.5 3.85 ;
      RECT 6.45 2.8 6.95 3.2 ;
      RECT 5.15 2.8 5.55 3.2 ;
      RECT 5.1 2.85 6.95 3.15 ;
      RECT 5.1 2.8 5.6 3.15 ;
      RECT 1.45 2.85 4.8 3.15 ;
      RECT 4.5 2.05 4.8 3.15 ;
      RECT 1.45 2.15 1.75 3.15 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 4.5 2.05 5.5 2.4 ;
      RECT 5 2 5.5 2.4 ;
    LAYER VIA12 ;
      RECT 6.57 2.87 6.83 3.13 ;
      RECT 5.22 2.87 5.48 3.13 ;
      RECT 5.12 2.07 5.38 2.33 ;
      RECT 3.37 3.57 3.63 3.83 ;
      RECT 1.47 2.22 1.73 2.48 ;
    LAYER MET1 ;
      RECT 5.45 3.5 5.75 5.2 ;
      RECT 4 3.5 6.15 3.8 ;
      RECT 5.85 1.55 6.15 3.8 ;
      RECT 4 2.75 4.3 3.8 ;
      RECT 3.85 2.75 4.3 3.2 ;
      RECT 5.45 1.55 6.15 1.8 ;
      RECT 5.45 0.95 5.75 1.8 ;
      RECT 3.45 3.5 3.75 5.2 ;
      RECT 3.15 1.55 3.45 3.9 ;
      RECT 3.45 0.95 3.75 1.8 ;
      RECT 1.45 0.95 1.75 5.2 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 6.45 2.85 6.95 3.15 ;
      RECT 5.1 2.8 5.6 3.25 ;
      RECT 5 2.05 5.5 2.35 ;
  END
END gf180mcu_osu_sc_gp9t3v3__lshifup
