# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_1 0 0 ;
  SIZE 3.2 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 3.2 6.35 ;
        RECT 1.4 3.6 1.75 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.2 0.7 ;
        RECT 1.4 0 1.75 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 2.95 1.55 3.25 ;
      LAYER Metal2 ;
        RECT 1.05 2.95 1.55 3.25 ;
        RECT 1.1 2.9 1.5 3.3 ;
      LAYER Via1 ;
        RECT 1.17 2.97 1.43 3.23 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 1.6 2.75 1.9 ;
        RECT 2.35 1.05 2.6 1.9 ;
        RECT 2.25 3.6 2.75 3.9 ;
        RECT 2.35 3.6 2.6 5.3 ;
      LAYER Metal2 ;
        RECT 2.25 3.55 2.75 3.95 ;
        RECT 2.25 1.55 2.75 1.95 ;
        RECT 2.35 1.55 2.65 3.95 ;
      LAYER Via1 ;
        RECT 2.37 3.62 2.63 3.88 ;
        RECT 2.37 1.62 2.63 1.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.55 1.05 0.8 5.3 ;
      RECT 0.55 2.25 2.2 2.55 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_1
