* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre = 0.0
.param sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_g5v0d10v5__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_g5v0d10v5 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__nfet_g5v0d10v5.0 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.995e-06 wmax = 1.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84203+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_0}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {107890+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_0}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_0}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_0}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_0}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_0}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_0}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_0}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_0}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_0}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_0}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_0+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_0}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_0}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_0}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_0}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_0}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_0}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_0}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_0}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_0}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.1 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.4995e-05 wmax = 1.5005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_1}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {97207+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_1}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_1}
+ ub = {2.0388e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_1}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_1}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_1}
+ a0 = {0.74065+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_1}
+ keta = {-0.027168+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_1}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_1}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_1}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_1}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_1+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_1}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_1}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33405+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_1}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 32.525
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_1}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_1}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_1}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_1}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_1}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.36273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_1}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4523e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.2 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.4995e-05 wmax = 1.5005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_2}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105660+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_2}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_2}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_2}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_2}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_2}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_2}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_2}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_2}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_2}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_2}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_2+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_2}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_2}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0792+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_2}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_2}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_2}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_2}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_2}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_2}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_2}
+ kt2 = -0.019151
+ at = 41664.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.3 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.85907+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019258+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_3}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {103150+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_3}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_3}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_3}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_3}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_3}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_3}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_3}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_3}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_3}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_3}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_3+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_3}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_3}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1563+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_3}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.7777e-5
+ alpha1 = 0.0
+ beta0 = 35.482
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_3}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_3}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_3}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_3}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_3}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_3}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.4 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83907+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019258+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_4}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {111130+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_4}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_4}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_4}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_4}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.041478+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_4}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_4}
+ keta = {-0.016843+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_4}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_4}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_4}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_4}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_4+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_4}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_4}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.43939+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_4}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.331e-5
+ alpha1 = 0.0
+ beta0 = 28.829
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_4}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_4}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_4}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_4}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_4}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_4}
+ kt2 = -0.019151
+ at = 20000.0
+ ute = -1.1947
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.5 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82471+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019258+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_5}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {116180+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_5}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_5}
+ ub = {1.7534e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_5}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_5}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.039819+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_5}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_5}
+ keta = {-0.025477+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_5}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_5}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_5}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_5}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_5+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_5}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_5}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.43939+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_5}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 26.7
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_5}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_5}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_5}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_5}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_5}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_5}
+ kt2 = -0.019151
+ at = 70000.0
+ ute = -1.1831
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.6 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.495e-06 wmax = 1.505e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.86603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_6}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {116860+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_6}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_6}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_6}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_6}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_6}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_6}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_6}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_6}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_6}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_6}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_6+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_6}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_6}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_6}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_6}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_6}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_6}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_6}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_6}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_6}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.7 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.85003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_7}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {107600+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_7}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_7}
+ ub = {1.4679e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_7}
+ uc = 4.6343e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_7}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.041406+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_7}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_7}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_7}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_7}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_7}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_7}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_7+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_7}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_7}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_7}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.8934e-5
+ alpha1 = 0.0
+ beta0 = 35.482
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_7}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_7}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_7}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_7}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_7}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_7}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.0908
+ ua1 = 3.0044e-9
+ ub1 = -3.3022e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.8 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.015173+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_8}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {110000+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_8}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_8}
+ ub = {1.5853e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_8}
+ uc = 6.5807e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_8}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.040476+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_8}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_8}
+ keta = {-0.021838+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_8}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_8}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_8}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_8}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_8+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_8}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_8}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_8}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.5046e-5
+ alpha1 = 0.0
+ beta0 = 29.568
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_8}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_8}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_8}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_8}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_8}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_8}
+ kt2 = -0.019151
+ at = 20000.0
+ ute = -1.1687
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.9 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.025187+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_9}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {111900+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_9}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_9}
+ ub = {1.617e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_9}
+ uc = 5.2646e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_9}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.038857+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_9}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_9}
+ keta = {-0.021838+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_9}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_9}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_9}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_9}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_9+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_9}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_9}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_9}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.1701e-5
+ alpha1 = 0.0
+ beta0 = 28.09
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_9}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_9}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_9}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_9}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_9}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_9}
+ kt2 = -0.019151
+ at = 40000.0
+ ute = -1.1687
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.10 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.025187+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_10}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {111900+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_10}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_10}
+ ub = {1.6817e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_10}
+ uc = 5.2646e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_10}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.038857+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_10}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_10}
+ keta = {-0.021838+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_10}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_10}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_10}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_10}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_10+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_10}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_10}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_10}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 3.0815e-5
+ alpha1 = 0.0
+ beta0 = 26.966
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_10}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_10}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_10}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_10}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_10}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_10}
+ kt2 = -0.019151
+ at = 150000.0
+ ute = -1.1687
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.11 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_11}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {118860+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_11}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_11}
+ ub = {1.5291e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_11}
+ uc = 4.6343e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_11}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_11}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_11}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_11}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_11}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_11}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_11}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_11+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_11}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_11}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_11}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_11}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_11}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_11}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_11}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_11}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_11}
+ kt2 = -0.019151
+ at = 40896.0
+ ute = -1.1428
+ ua1 = 3.0044e-9
+ ub1 = -1.7594e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.12 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.86947+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019258+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_12}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109350+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_12}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_12}
+ ub = {1.5291e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_12}
+ uc = 5.9319e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_12}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_12}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_12}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_12}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_12}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_12}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_12}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_12+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_12}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_12}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.7473+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_12}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.9675e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_12}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_12}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_12}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_12}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_12}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_12}
+ kt2 = -0.019151
+ at = 38400.0
+ ute = -1.2991
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.13 nmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 9.95e-07 wmax = 1.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.015173+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_13}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {111900+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_13}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_13}
+ ub = {1.4679e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_13}
+ uc = 6.5807e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_13}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.042162+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_13}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_13}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_13}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_13}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_13}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_13}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_13+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_13}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_13}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_13}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 3.2414e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_13}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_13}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_13}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_13}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_13}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_13}
+ kt2 = -0.019151
+ at = 29000.0
+ ute = -1.2471
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.14 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 1.9995e-05 wmax = 2.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_14}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {94207+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_14}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_14}
+ ub = {2.0388e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_14}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_14}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_14}
+ a0 = {0.74065+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_14}
+ keta = {-0.027168+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_14}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_14}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_14}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_14}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_14+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_14}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_14}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33405+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_14}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 32.5
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_14}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_14}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_14}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_14}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_14}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.36273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_14}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4523e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.15 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 1.9995e-05 wmax = 2.0005e-5
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_15}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105660+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_15}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_15}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_15}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_15}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_15}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_15}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_15}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_15}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_15}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_15}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_15+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_15}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_15}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_15}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_15}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_15}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_15}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_15}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_15}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_15}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4025e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.16 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.018091+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_16}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {101100+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_16}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_16}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_16}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_16}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_16}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_16}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_16}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_16}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_16}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_16}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_16+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_16}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_16}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.89936+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_16}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.8807e-5
+ alpha1 = 0.0
+ beta0 = 34.003
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_16}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_16}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_16}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_16}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_16}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_16}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.17 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.018091+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_17}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100100+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_17}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_17}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_17}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_17}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.042006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_17}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_17}
+ keta = {-0.03033+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_17}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_17}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_17}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_17}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_17+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_17}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_17}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.89936+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_17}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 29.9
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_17}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_17}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_17}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_17}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_17}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_17}
+ kt2 = -0.019151
+ at = 10000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.18 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.018091+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_18}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {86056+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_18}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_18}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_18}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_18}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.0414+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_18}
+ a0 = {0.96509+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_18}
+ keta = {-0.03033+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_18}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_18}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_18}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_18}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_18+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_18}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_18}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.89936+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_18}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.3888e-5
+ alpha1 = 0.0
+ beta0 = 26.7
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_18}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_18}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_18}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_18}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_18}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_18}
+ kt2 = -0.019151
+ at = 60000.0
+ ute = -1.2586
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.19 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.018091+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_19}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {78024+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_19}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_19}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_19}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_19}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.0414+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_19}
+ a0 = {0.96509+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_19}
+ keta = {-0.03033+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_19}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_19}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_19}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_19}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_19+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_19}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_19}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.89936+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_19}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 23.8
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_19}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_19}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_19}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_19}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_19}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.40273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_19}
+ kt2 = -0.019151
+ at = 113600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.20 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83803+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_20}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {109890+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_20}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_20}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_20}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_20}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_20}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_20}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_20}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_20}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_20}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_20}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_20+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_20}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_20}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_20}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_20}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_20}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_20}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_20}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_20}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_20}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.5525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.21 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 2.995e-06 wmax = 3.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84203+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.020425+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_21}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105490+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_21}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_21}
+ ub = {1.8689e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_21}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_21}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_21}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_21}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_21}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_21}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_21}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_21}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_21+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_21}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_21}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_21}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.8228e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_21}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_21}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_21}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_21}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_21}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_21}
+ kt2 = -0.019151
+ at = 38400.0
+ ute = -1.2991
+ ua1 = 2.0117e-9
+ ub1 = -1.513e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.22 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_22}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {97207+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_22}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_22}
+ ub = {1.8265e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_22}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_22}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_22}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_22}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_22}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_22}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_22}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_22}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_22+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_22}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_22}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.89936+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_22}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.8934e-5
+ alpha1 = 0.0
+ beta0 = 35.6
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_22}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_22}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_22}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_22}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_22}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_22}
+ kt2 = -0.019151
+ at = 30000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.23 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82703+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_23}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {103550+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_23}
+ ua = {3.3055e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_23}
+ ub = {1.7534e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_23}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_23}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044934+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_23}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_23}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_23}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_23}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_23}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_23}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_23+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_23}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_23}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2052+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_23}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 29.568
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_23}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_23}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_23}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_23}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_23}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_23}
+ kt2 = -0.019151
+ at = 20000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.24 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82903+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_24}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {102820+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_24}
+ ua = {6.611e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_24}
+ ub = {1.8235e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_24}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_24}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044934+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_24}
+ a0 = {0.83043+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_24}
+ keta = {-0.023051+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_24}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.14102+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_24}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_24}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_24}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_24+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_24}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_24}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2052+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_24}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.5624e-5
+ alpha1 = 0.0
+ beta0 = 26.611
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_24}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_24}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_24}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_24}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_24}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_24}
+ kt2 = -0.019151
+ at = 80000.0
+ ute = -1.2586
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.25 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.8206+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_25}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100190+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_25}
+ ua = {6.611e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_25}
+ ub = {1.8235e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_25}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_25}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044934+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_25}
+ a0 = {0.83043+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_25}
+ keta = {-0.023051+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_25}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.13538+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_25}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_25}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_25}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_25+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_25}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_25}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.2052+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_25}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.0706e-5
+ alpha1 = 0.0
+ beta0 = 22.915
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_25}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_25}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_25}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_25}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_25}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.40273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_25}
+ kt2 = -0.019151
+ at = 152000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.26 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84303+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_26}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108890+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_26}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_26}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_26}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_26}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_26}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_26}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_26}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_26}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_26}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_26}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_26+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_26}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_26}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_26}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_26}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_26}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_26}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_26}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_26}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_26}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.5525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.27 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_27}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105140+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_27}
+ ua = {-8.3888e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_27}
+ ub = {1.7534e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_27}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_27}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044934+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_27}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_27}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_27}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_27}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_27}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_27}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_27+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_27}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_27}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.026+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_27}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.765e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_27}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_27}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_27}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_27}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_27}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_27}
+ kt2 = -0.019151
+ at = 38400.0
+ ute = -1.2991
+ ua1 = 2.0117e-9
+ ub1 = -1.347e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.28 nmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 4.995e-06 wmax = 5.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_28}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {101100+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_28}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_28}
+ ub = {1.7534e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_28}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_28}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_28}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_28}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_28}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_28}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_28}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_28}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_28+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_28}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_28}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.82741+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_28}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.0254e-5
+ alpha1 = 0.0
+ beta0 = 35.482
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_28}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_28}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_28}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_28}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_28}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_28}
+ kt2 = -0.019151
+ at = 29000.0
+ ute = -1.2471
+ ua1 = 2.0117e-9
+ ub1 = -1.257e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.29 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_29}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {101430+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_29}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_29}
+ ub = {2.0388e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_29}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_29}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_29}
+ a0 = {1.2569+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_29}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_29}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_29}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_29}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_29}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_29+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_29}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_29}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.71949+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_29}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.331e-5
+ alpha1 = 0.0
+ beta0 = 32.8
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_29}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_29}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_29}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_29}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_29}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_29}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.30 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82403+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_30}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {108110+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_30}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_30}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_30}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_30}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_30}
+ a0 = {1.2569+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_30}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_30}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_30}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_30}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_30}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_30+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_30}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_30}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.20557+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_30}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 29.568
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_30}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_30}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_30}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_30}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_30}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_30}
+ kt2 = -0.019151
+ at = 16000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.31 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.82603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_31}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100660+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_31}
+ ua = {-1.7976e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_31}
+ ub = {1.9964e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_31}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_31}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_31}
+ a0 = {0.85287+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_31}
+ keta = {-0.025533+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_31}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.14102+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_31}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_31}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_31}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_31+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_31}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_31}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.41114+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_31}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 26.6
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_31}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_31}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_31}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_31}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_31}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_31}
+ kt2 = -0.019151
+ at = 80000.0
+ ute = -1.2586
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.32 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.81703+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_32}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105660+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_32}
+ ua = {-6.2916e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_32}
+ ub = {2.0813e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_32}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_32}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_32}
+ a0 = {0.94535+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_32}
+ keta = {-0.02132+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_32}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.14743+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_32}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_32}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_32}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_32+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_32}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_32}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.33405+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_32}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 24.0
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_32}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_32}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_32}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_32}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_32}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.40273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_32}
+ kt2 = -0.019151
+ at = 160000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.33 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_33}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {105660+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_33}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_33}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_33}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_33}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_33}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_33}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_33}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_33}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_33}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_33}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_33+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_33}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_33}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_33}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_33}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_33}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_33}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_33}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_33}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_33}
+ kt2 = -0.019151
+ at = 40000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.5525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.34 nmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 6.995e-06 wmax = 7.005e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.029179+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_34}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {100430+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_34}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_34}
+ ub = {2.1238e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_34}
+ uc = 6.6204e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_34}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_34}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_34}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_34}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_34}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_34}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_34}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_34+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_34}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_34}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.0278+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_34}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.736e-5
+ alpha1 = 0.0
+ beta0 = 35.482
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_34}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_34}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_34}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_34}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_34}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_34}
+ kt2 = -0.019151
+ at = 29000.0
+ ute = -1.2471
+ ua1 = 2.0117e-9
+ ub1 = -1.447e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.35 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.844+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.016501+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_35}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {123750+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_35}
+ ua = {-7.49e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_35}
+ ub = {1.5903e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_35}
+ uc = 6.0802e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_35}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.048606+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_35}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_35}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_35}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_35}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_35}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_35}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_35+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_35}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_35}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1363+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_35}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 32.525
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_35}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_35}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_35}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_35}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_35}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_35}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.36 nmos
* DC IV MOS Parameters
+ lmin = 1.9995e-05 lmax = 2.0005e-05 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.835+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.031405+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_36}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {128700+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_36}
+ ua = {0+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_36}
+ ub = {1.9579e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_36}
+ uc = 7.8119e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_36}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044796+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_36}
+ a0 = {1.104+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_36}
+ keta = {-0.01489+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_36}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_36}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_36}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_36}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_36+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_36}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_36}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.49997+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_36}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 3.7422e-5
+ alpha1 = 0.0
+ beta0 = 24.268
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_36}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_36}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_36}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_36}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_36}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.38773+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_36}
+ kt2 = -0.019151
+ at = 260000.0
+ ute = -1.0389
+ ua1 = 3.0044e-9
+ ub1 = -3.4523e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.37 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.025742+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_37}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {120700+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_37}
+ ua = {-7.49e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_37}
+ ub = {1.8129e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_37}
+ uc = 6.0802e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_37}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.046662+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_37}
+ a0 = {0.80798+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_37}
+ keta = {-0.02068+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_37}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_37}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_37}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_37}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_37+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_37}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_37}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.49997+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_37}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.5914e-5
+ alpha1 = 0.0
+ beta0 = 29.923
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_37}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_37}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_37}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_37}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_37}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_37}
+ kt2 = -0.019151
+ at = 20000.0
+ ute = -1.1687
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.38 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.838+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_38+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.031405+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_38}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {122700+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_38}
+ ua = {0+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_38}
+ ub = {1.8129e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_38}
+ uc = 5.3506e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_38}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044796+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_38}
+ a0 = {0.90494+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_38}
+ keta = {-0.02068+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_38}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_38}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_38}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_38}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_38+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_38+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_38}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_38}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.49997+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_38}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4641e-5
+ alpha1 = 0.0
+ beta0 = 26.332
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_38}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_38}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_38}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_38}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_38}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_38}
+ kt2 = -0.019151
+ at = 80000.0
+ ute = -1.1327
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.39 nmos
* DC IV MOS Parameters
+ lmin = 7.995e-06 lmax = 8.005e-06 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.843+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_39+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.031405+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_39}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {128700+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_39}
+ ua = {0+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_39}
+ ub = {1.9579e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_39}
+ uc = 7.8119e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_39}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044796+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_39}
+ a0 = {0.90494+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_39}
+ keta = {-0.01489+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_39}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_39}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_39}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_39}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_39+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_39+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_39}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_39}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.49997+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_39}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.079e-5
+ alpha1 = 0.0
+ beta0 = 25.279
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_39}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_39}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_39}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_39}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_39}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.40273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_39}
+ kt2 = -0.019151
+ at = 192000.0
+ ute = -1.1168
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.40 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.804+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_40+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.013096+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_40}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {132070+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_40}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_40}
+ ub = {1.5903e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_40}
+ uc = 3.8001e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_40}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.048606+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_40}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_40}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_40}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_40}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_40}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_40}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_40+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_40+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_40}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_40}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.7216+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_40}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_40}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_40}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_40}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_40}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_40}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.33573+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_40}
+ kt2 = -0.019151
+ at = 49600.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.41 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84464+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_41+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.0072604+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_41}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {125700+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_41}
+ ua = {-9.8868e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_41}
+ ub = {1.4758e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_41}
+ uc = 5.229e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_41}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.049906+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_41}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_41}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_41}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_41}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_41}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_41}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_41+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_41+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_41}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_41}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.5681+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_41}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 9.8376e-6
+ alpha1 = 0.0
+ beta0 = 33.826
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_41}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_41}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_41}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_41}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_41}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_41}
+ kt2 = -0.019151
+ at = 38400.0
+ ute = -1.2991
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.42 nmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 4.15e-07 wmax = 4.25e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.870+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_42+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.0072604+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_42}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {123750+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_42}
+ ua = {-9.8868e-011+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_42}
+ ub = {1.2722e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_42}
+ uc = 5.229e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_42}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.048606+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_42}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_42}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_42}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_42}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_42}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_42}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_42+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_42+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_42}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_42}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1363+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_42}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 9.8376e-6
+ alpha1 = 0.0
+ beta0 = 32.525
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_42}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_42}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_42}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_42}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_42}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_42}
+ kt2 = -0.019151
+ at = 29000.0
+ ute = -1.2471
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.43 nmos
* DC IV MOS Parameters
+ lmin = 9.95e-07 lmax = 1.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_43+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019842+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_43}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {106500+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_43}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_43}
+ ub = {1.5291e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_43}
+ uc = 5.7002e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_43}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_43}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_43}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_43}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_43}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_43}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_43}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_43+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_43+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_43}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_43}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_43}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.8066e-5
+ alpha1 = 0.0
+ beta0 = 35.482
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_43}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_43}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_43}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_43}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_43}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_43}
+ kt2 = -0.019151
+ at = 24000.0
+ ute = -1.2986
+ ua1 = 3.0044e-9
+ ub1 = -3.4525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.81e-6
+ sbref = 2.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.44 nmos
* DC IV MOS Parameters
+ lmin = 1.995e-06 lmax = 2.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.85803+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_44+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.023414+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_44}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {111000+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_44}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_44}
+ ub = {1.6514e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_44}
+ uc = 5.7002e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_44}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.041478+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_44}
+ a0 = {0.67332+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_44}
+ keta = {-0.020254+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_44}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_44}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_44}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_44}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_44+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_44+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_44}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_44}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.20557+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_44}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.8066e-5
+ alpha1 = 0.0
+ beta0 = 31.224
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_44}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_44}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_44}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_44}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_44}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37273+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_44}
+ kt2 = -0.019151
+ at = 20000.0
+ ute = -1.1687
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.45 nmos
* DC IV MOS Parameters
+ lmin = 3.995e-06 lmax = 4.005e-06 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_45+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.023414+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_45}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {101000+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_45}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_45}
+ ub = {1.7175e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_45}
+ uc = 5.7002e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_45}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.039819+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_45}
+ a0 = {0.80798+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_45}
+ keta = {-0.020254+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_45}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_45}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_45}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_45}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_45+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_45+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_45}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_45}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {0.20557+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_45}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 2.8066e-5
+ alpha1 = 0.0
+ beta0 = 28.726
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_45}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_45}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_45}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_45}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_45}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.39073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_45}
+ kt2 = -0.019151
+ at = 60000.0
+ ute = -1.1327
+ ua1 = 3.0044e-9
+ ub1 = -3.7525e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.46 nmos
* DC IV MOS Parameters
+ lmin = 4.95e-07 lmax = 5.05e-07 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope1/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.84003+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_46+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019842+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_46}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {121610+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_46}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_46}
+ ub = {1.5291e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_46}
+ uc = 3.8001e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_46}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.045006+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_46}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_46}
+ keta = {-0.01066+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_46}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_46}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_46}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_46}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_46+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_46+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_46}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_46}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.2848+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_46}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.4467e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_46}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_46}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_46}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_46}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_46}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.35073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_46}
+ kt2 = -0.019151
+ at = 40896.0
+ ute = -1.1428
+ ua1 = 3.0044e-9
+ ub1 = -1.9993e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 1.81e-6
+ sbref = 1.81e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.47 nmos
* DC IV MOS Parameters
+ lmin = 7.95e-07 lmax = 8.05e-07 wmin = 7.45e-07 wmax = 7.55e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.83603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_47+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019842+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_47}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {116750+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_47}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_47}
+ ub = {1.5903e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_47}
+ uc = 6.0042e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_47}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.043206+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_47}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_47}
+ keta = {-0.0044772+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_47}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_47}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_47}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_47}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_47+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_47+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_47}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_47}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1049+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_47}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 3.2296e-5
+ alpha1 = 0.0
+ beta0 = 36.96
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_47}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_47}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_47}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_47}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_47}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_47}
+ kt2 = -0.019151
+ at = 29000.0
+ ute = -1.2471
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.41e-6
+ sbref = 2.41e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__nfet_g5v0d10v5.48 nmos
* DC IV MOS Parameters
+ lmin = 5.95e-07 lmax = 6.05e-07 wmin = 6.95e-07 wmax = 7.05e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 1.16e-8
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = {7.6507e-008+sky130_fd_pr__nfet_g5v0d10v5__lint_diff}
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = {2.1346e-008+sky130_fd_pr__nfet_g5v0d10v5__wint_diff}
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -4.1292e-9
+ dwb = -1.6944e-9
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.794
+ rnoib = 0.38
+ tnoia = 7.50e+6
+ tnoib = 7.2e+6
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {1.16e-008*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult+MC_MM_SWITCH*(1.16e-08*sky130_fd_pr__nfet_g5v0d10v5__toxe_mult*(sky130_fd_pr__nfet_g5v0d10v5__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = {1*sky130_fd_pr__nfet_g5v0d10v5__rshn_mult}
* Threshold Voltage Parameters
+ vth0 = {0.85603+sky130_fd_pr__nfet_g5v0d10v5__vth0_diff_48+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__vth0_slope/sqrt(1))}
+ k1 = 0.88325
+ k2 = {-0.019842+sky130_fd_pr__nfet_g5v0d10v5__k2_diff_48}
+ k3 = -0.884
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.19251
+ dvt0w = 0.16
+ dvt1w = 6909100.0
+ dvt2w = -0.036016
+ w0 = 0.0
+ k3b = 0.43
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 2.5e-8
+ lpeb = -2.182e-7
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = {123420+sky130_fd_pr__nfet_g5v0d10v5__vsat_diff_48}
+ ua = {-1.498e-010+sky130_fd_pr__nfet_g5v0d10v5__ua_diff_48}
+ ub = {1.7175e-018+sky130_fd_pr__nfet_g5v0d10v5__ub_diff_48}
+ uc = 6.4845e-11
+ rdsw = {724.62+sky130_fd_pr__nfet_g5v0d10v5__rdsw_diff_48}
+ prwb = 0.05626
+ prwg = 0.048
+ wr = 1.0
+ u0 = {0.044934+sky130_fd_pr__nfet_g5v0d10v5__u0_diff_48}
+ a0 = {1.1222+sky130_fd_pr__nfet_g5v0d10v5__a0_diff_48}
+ keta = {-0.0044772+sky130_fd_pr__nfet_g5v0d10v5__keta_diff_48}
+ a1 = 0.0
+ a2 = 0.65972622
+ ags = {0.16025+sky130_fd_pr__nfet_g5v0d10v5__ags_diff_48}
+ b0 = {3.2933e-008+sky130_fd_pr__nfet_g5v0d10v5__b0_diff_48}
+ b1 = {0+sky130_fd_pr__nfet_g5v0d10v5__b1_diff_48}
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.20613+sky130_fd_pr__nfet_g5v0d10v5__voff_diff_48+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__voff_slope/sqrt(1))}
+ nfactor = {0.5412+sky130_fd_pr__nfet_g5v0d10v5__nfactor_diff_48+MC_MM_SWITCH*(sky130_fd_pr__nfet_g5v0d10v5__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = {0+sky130_fd_pr__nfet_g5v0d10v5__tvoff_diff_48}
+ cit = -0.0008
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0
+ eta0 = {0.032+sky130_fd_pr__nfet_g5v0d10v5__eta0_diff_48}
+ etab = -0.01932
+ dsub = 0.504
* BSIM4 - Sub-threshold parameters
+ voffl = -4.2579486e-7
+ minv = 0.0
* Rout Parameters
+ pclm = {1.1049+sky130_fd_pr__nfet_g5v0d10v5__pclm_diff_48}
+ pdiblc1 = 0.21098
+ pdiblc2 = 0.0002
+ pdiblcb = -0.26831
+ drout = 0.36075
+ pscbe1 = 9.3731e+8
+ pscbe2 = 1.68e-6
+ pvag = 1.99
+ delta = 0.0246
+ alpha0 = 1.9378e-5
+ alpha1 = 0.0
+ beta0 = 36.6
* BSIM4 - Rout Parameters
+ fprout = 10.125
+ pdits = {0+sky130_fd_pr__nfet_g5v0d10v5__pdits_diff_48}
+ pditsl = 0.0
+ pditsd = {0+sky130_fd_pr__nfet_g5v0d10v5__pditsd_diff_48}
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = {5.06e-011+sky130_fd_pr__nfet_g5v0d10v5__agidl_diff_48}
+ bgidl = {1.058e009+sky130_fd_pr__nfet_g5v0d10v5__bgidl_diff_48}
+ cgidl = {4000+sky130_fd_pr__nfet_g5v0d10v5__cgidl_diff_48}
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 1.16e-8
* Temperature Effects Parameters
+ kt1 = {-0.37073+sky130_fd_pr__nfet_g5v0d10v5__kt1_diff_48}
+ kt2 = -0.019151
+ at = 38400.0
+ ute = -1.2991
+ ua1 = 2.0117e-9
+ ub1 = -1.8012e-18
+ uc1 = -5.9821e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 2.6e+41
+ noib = 0.0
+ noic = 0.0
+ em = 4.1000000e+7
+ af = 1.0
+ ef = 0.89
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.0773
+ jss = 0.000375
+ jsws = 5.84e-11
+ xtis = 0.76
+ bvs = 12.636
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001344
+ tpbsw = 0.00099005
+ tpbswg = 0.0
+ tcj = 0.00067434
+ tcjsw = 0.0002493
+ tcjswg = 0.0
+ cgdo = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgso = {3.0674e-010*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgbo = 0.0
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cgdl = {5e-011*sky130_fd_pr__nfet_g5v0d10v5__overlap_mult}
+ cf = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ dlc = {6.5995e-008+sky130_fd_pr__nfet_g5v0d10v5__dlc_diff+sky130_fd_pr__nfet_g5v0d10v5__dlc_rotweak}
+ dwc = {0+sky130_fd_pr__nfet_g5v0d10v5__dwc_diff}
+ vfbcv = -1.0
+ acde = 0.4176
+ moin = 15.0
+ noff = 4.0
+ voffcv = -0.4104
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = {0.0008512*sky130_fd_pr__nfet_g5v0d10v5__ajunction_mult}
+ mjs = 0.295
+ pbs = 0.72468
+ cjsws = {8.5204e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjsws = 0.037586
+ pbsws = 0.29067
+ cjswgs = {5.4e-011*sky130_fd_pr__nfet_g5v0d10v5__pjunction_mult}
+ mjswgs = 0.78692
+ pbswgs = 0.54958
* Stress Parameters
+ saref = 2.02e-6
+ sbref = 2.01e-6
+ wlod = {0+sky130_fd_pr__nfet_g5v0d10v5__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__ku0_diff}
+ lku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__lku0_diff}
+ wku0 = {0+sky130_fd_pr__nfet_g5v0d10v5__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__nfet_g5v0d10v5__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__nfet_g5v0d10v5
