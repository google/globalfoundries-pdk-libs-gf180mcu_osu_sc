VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addf_1 0 0 ;
  SIZE 14 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 14 6.15 ;
        RECT 12.35 4.7 12.6 6.15 ;
        RECT 10.75 4.7 11 6.15 ;
        RECT 6.5 4.7 6.75 6.15 ;
        RECT 4.8 4.7 5.05 6.15 ;
        RECT 1.4 4.7 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14 0.6 ;
        RECT 12.35 0 12.6 1.4 ;
        RECT 10.75 0 11 1.4 ;
        RECT 6.5 0 6.75 1.4 ;
        RECT 4.8 0 5.05 1.4 ;
        RECT 1.4 0 1.65 1.4 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.7 2.35 9.2 2.65 ;
        RECT 6.4 3.05 9.1 3.35 ;
        RECT 8.8 2.35 9.1 3.35 ;
        RECT 6.4 2.35 6.7 3.35 ;
        RECT 3.2 2.35 6.7 2.65 ;
        RECT 2.15 3.1 3.45 3.4 ;
        RECT 3.2 2.35 3.45 3.4 ;
        RECT 2.15 2.2 2.4 3.4 ;
        RECT 0.6 2.2 2.4 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.85 3.6 9.95 3.9 ;
        RECT 9.65 2.9 9.95 3.9 ;
        RECT 5.85 2.9 6.15 3.9 ;
        RECT 3.7 3 6.15 3.3 ;
        RECT 1.6 3.65 4 3.95 ;
        RECT 3.7 2.9 4 3.95 ;
        RECT 1.6 2.75 1.9 3.95 ;
      LAYER MET2 ;
        RECT 1.5 2.85 2 3.15 ;
        RECT 1.55 2.8 1.95 3.2 ;
      LAYER VIA12 ;
        RECT 1.62 2.87 1.88 3.13 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.75 2.25 10.6 2.55 ;
        RECT 9.75 1.8 10.05 2.55 ;
        RECT 2.65 1.8 10.05 2.1 ;
        RECT 7.05 1.8 7.35 2.75 ;
        RECT 2.65 1.8 2.95 2.6 ;
      LAYER MET2 ;
        RECT 2.55 2.2 3.05 2.5 ;
        RECT 2.6 2.15 3 2.55 ;
      LAYER VIA12 ;
        RECT 2.67 2.22 2.93 2.48 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.2 3 13.75 3.3 ;
        RECT 13.2 2.95 13.65 3.35 ;
        RECT 13.2 0.95 13.45 5.2 ;
      LAYER MET2 ;
        RECT 13.25 3 13.75 3.3 ;
        RECT 13.3 2.95 13.7 3.35 ;
      LAYER VIA12 ;
        RECT 13.37 3.02 13.63 3.28 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.6 3 12.05 3.3 ;
        RECT 11.6 2.95 11.9 3.35 ;
        RECT 11.6 0.95 11.85 5.2 ;
      LAYER MET2 ;
        RECT 11.55 3 12.05 3.3 ;
        RECT 11.6 2.95 12 3.35 ;
      LAYER VIA12 ;
        RECT 11.67 3.02 11.93 3.28 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 3.1 4.75 3.4 5.2 ;
      RECT 3.05 4.75 3.45 5.15 ;
      RECT 3 4.8 12.85 5.1 ;
      RECT 12.55 2.25 12.85 5.1 ;
      RECT 3.75 1.05 4.05 5.1 ;
      RECT 12.5 2.3 12.9 2.7 ;
      RECT 7.85 2.3 8.25 2.7 ;
      RECT 12.45 2.35 12.95 2.65 ;
      RECT 3.75 2.35 8.3 2.65 ;
      RECT 3.1 0.95 3.4 1.45 ;
      RECT 3.05 1 3.45 1.4 ;
      RECT 3.05 1.05 4.05 1.35 ;
      RECT 8.15 4.1 8.55 4.5 ;
      RECT 8.1 4.15 11.25 4.45 ;
      RECT 10.95 2.25 11.25 4.45 ;
      RECT 8.85 1.05 9.15 4.45 ;
      RECT 10.9 2.3 11.3 2.7 ;
      RECT 8.15 1 8.55 1.4 ;
      RECT 8.1 1.05 9.15 1.35 ;
      RECT 7.3 0.95 7.6 1.45 ;
      RECT 5.65 0.95 5.95 1.45 ;
      RECT 7.25 1 7.65 1.4 ;
      RECT 5.6 1 6 1.4 ;
      RECT 5.6 1.05 7.65 1.35 ;
      RECT 2.2 0.95 2.5 1.45 ;
      RECT 0.5 0.95 0.8 1.45 ;
      RECT 2.15 1 2.55 1.4 ;
      RECT 0.45 1 0.85 1.4 ;
      RECT 0.45 1.05 2.55 1.35 ;
    LAYER VIA12 ;
      RECT 12.57 2.37 12.83 2.63 ;
      RECT 10.97 2.37 11.23 2.63 ;
      RECT 8.22 1.07 8.48 1.33 ;
      RECT 8.22 4.17 8.48 4.43 ;
      RECT 7.92 2.37 8.18 2.63 ;
      RECT 7.32 1.07 7.58 1.33 ;
      RECT 5.67 1.07 5.93 1.33 ;
      RECT 3.12 1.07 3.38 1.33 ;
      RECT 3.12 4.82 3.38 5.08 ;
      RECT 2.22 1.07 2.48 1.33 ;
      RECT 0.52 1.07 0.78 1.33 ;
    LAYER MET1 ;
      RECT 7.35 4.2 7.6 5.2 ;
      RECT 5.65 4.2 5.9 5.2 ;
      RECT 5.65 4.2 7.6 4.45 ;
      RECT 2.25 4.2 2.5 5.2 ;
      RECT 0.55 4.2 0.8 5.2 ;
      RECT 0.55 4.2 2.5 4.45 ;
      RECT 12.45 2.35 12.95 2.65 ;
      RECT 10.85 2.35 11.35 2.65 ;
      RECT 8.1 4.15 8.6 4.45 ;
      RECT 8.2 0.95 8.5 1.45 ;
      RECT 7.8 2.35 8.3 2.65 ;
      RECT 7.3 0.95 7.6 1.45 ;
      RECT 5.65 0.95 5.95 1.45 ;
      RECT 3.1 0.95 3.4 1.45 ;
      RECT 3.1 4.7 3.4 5.2 ;
      RECT 2.2 0.95 2.5 1.45 ;
      RECT 0.5 0.95 0.8 1.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addf_1

MACRO gf180mcu_osu_sc_gp9t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addh_1 0 0 ;
  SIZE 8.6 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.6 6.15 ;
        RECT 6.65 4.5 6.9 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.6 0.6 ;
        RECT 6.65 0 6.9 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 2.2 4.4 2.5 ;
        RECT 1.5 2.2 2 2.5 ;
      LAYER MET2 ;
        RECT 3.9 2.15 4.4 2.55 ;
        RECT 1.5 2.2 4.4 2.5 ;
        RECT 1.5 2.15 2 2.55 ;
      LAYER VIA12 ;
        RECT 1.62 2.22 1.88 2.48 ;
        RECT 4.02 2.22 4.28 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 1.9 5.5 2.4 ;
        RECT 2.35 2.15 2.85 2.45 ;
        RECT 2.35 1.55 2.85 1.85 ;
        RECT 2.45 1.55 2.75 2.45 ;
      LAYER MET2 ;
        RECT 5.15 1.95 5.55 2.35 ;
        RECT 5.2 1.55 5.5 2.4 ;
        RECT 5.15 1.55 5.5 2.35 ;
        RECT 2.35 1.55 5.5 1.85 ;
        RECT 2.4 1.5 2.8 1.9 ;
      LAYER VIA12 ;
        RECT 2.47 1.57 2.73 1.83 ;
        RECT 5.22 2.02 5.48 2.28 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
        RECT 0.55 0.95 0.8 5.2 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.7 2.85 8.2 3.15 ;
        RECT 7.75 2.8 8.1 3.2 ;
        RECT 7.5 3.5 8 5.2 ;
        RECT 7.75 0.95 8 5.2 ;
      LAYER MET2 ;
        RECT 7.7 2.8 8.2 3.2 ;
      LAYER VIA12 ;
        RECT 7.82 2.87 8.08 3.13 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 6.3 2.95 6.8 3.35 ;
      RECT 3 2.9 3.5 3.3 ;
      RECT 3 2.95 6.8 3.25 ;
    LAYER VIA12 ;
      RECT 6.42 3.02 6.68 3.28 ;
      RECT 3.12 2.97 3.38 3.23 ;
    LAYER MET1 ;
      RECT 5.55 3.5 6.05 5.2 ;
      RECT 5.55 2.75 5.8 5.2 ;
      RECT 4.7 2.75 6.05 3 ;
      RECT 5.75 2.5 6.75 2.75 ;
      RECT 4.7 1.35 4.95 3 ;
      RECT 6.5 2.2 7.25 2.5 ;
      RECT 5.55 0.85 5.8 1.45 ;
      RECT 3.85 0.85 4.1 1.45 ;
      RECT 3.85 0.85 5.8 1.1 ;
      RECT 2.25 2.95 2.5 5.2 ;
      RECT 1.05 2.95 3.5 3.25 ;
      RECT 3.1 0.95 3.35 3.25 ;
      RECT 6.3 3 6.8 3.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addh_1

MACRO gf180mcu_osu_sc_gp9t3v3__and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__and2_1 0 0 ;
  SIZE 4.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.1 6.15 ;
        RECT 2.25 3.5 2.7 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.1 0.6 ;
        RECT 2.1 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.2 1.1 2.5 ;
        RECT 0.65 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.8 2.45 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 3.5 3.8 3.8 ;
        RECT 3.3 3.45 3.7 3.85 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 3.3 3.45 3.8 3.85 ;
      LAYER VIA12 ;
        RECT 3.42 3.52 3.68 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.45 1.65 5.2 ;
      RECT 2.75 2.1 3.05 2.6 ;
      RECT 1.4 2.2 3.05 2.5 ;
      RECT 0.7 1.45 1.65 1.7 ;
      RECT 0.7 0.95 0.95 1.7 ;
  END
END gf180mcu_osu_sc_gp9t3v3__and2_1

MACRO gf180mcu_osu_sc_gp9t3v3__aoi21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi21_1 0 0 ;
  SIZE 3.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.9 6.15 ;
        RECT 1.4 4.25 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.95 0 3.2 1.4 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 2.2 2.85 2.5 ;
      LAYER MET2 ;
        RECT 2.35 2.15 2.85 2.55 ;
      LAYER VIA12 ;
        RECT 2.47 2.22 2.73 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 3.5 3.5 3.8 ;
        RECT 3.1 1.65 3.35 5.2 ;
        RECT 2.1 1.65 3.35 1.9 ;
        RECT 2.1 0.95 2.35 1.9 ;
      LAYER MET2 ;
        RECT 3 3.45 3.5 3.85 ;
      LAYER VIA12 ;
        RECT 3.12 3.52 3.38 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.25 3.75 2.5 5.2 ;
      RECT 0.55 3.75 0.8 5.2 ;
      RECT 0.55 3.75 2.5 4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi21_1

MACRO gf180mcu_osu_sc_gp9t3v3__aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi22_1 0 0 ;
  SIZE 5.4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.4 6.15 ;
        RECT 1.4 4.25 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.4 0.6 ;
        RECT 3.5 0 3.75 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.4 2.85 2.9 3.15 ;
      LAYER MET2 ;
        RECT 2.4 2.8 2.9 3.2 ;
      LAYER VIA12 ;
        RECT 2.52 2.87 2.78 3.13 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 2.85 3.8 3.15 ;
      LAYER MET2 ;
        RECT 3.3 2.8 3.8 3.2 ;
      LAYER VIA12 ;
        RECT 3.42 2.87 3.68 3.13 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.5 4.05 4.8 4.55 ;
        RECT 4.55 2.05 4.8 4.55 ;
        RECT 2.1 2.05 4.8 2.3 ;
        RECT 2.1 0.95 2.35 2.3 ;
        RECT 3 4.15 3.5 4.45 ;
        RECT 3.1 4.15 3.35 5.2 ;
      LAYER MET2 ;
        RECT 4.45 4.05 4.85 4.55 ;
        RECT 3 4.15 4.85 4.45 ;
        RECT 3 4.1 3.5 4.5 ;
      LAYER VIA12 ;
        RECT 3.12 4.17 3.38 4.43 ;
        RECT 4.52 4.17 4.78 4.43 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.95 3.65 4.25 5.2 ;
      RECT 2.25 3.65 2.5 5.2 ;
      RECT 0.55 3.65 0.8 5.2 ;
      RECT 0.55 3.65 4.25 3.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi22_1

MACRO gf180mcu_osu_sc_gp9t3v3__aoi31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi31_1 0 0 ;
  SIZE 4.95 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.95 6.15 ;
        RECT 2.25 4.25 2.5 6.15 ;
        RECT 0.55 3.75 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.95 0.6 ;
        RECT 3.8 0 4.05 1.8 ;
        RECT 0.95 0 1.2 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 2.85 3 3.15 ;
      LAYER MET2 ;
        RECT 2.5 2.8 3 3.2 ;
      LAYER VIA12 ;
        RECT 2.62 2.87 2.88 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 2.85 1.25 3.15 ;
      LAYER MET2 ;
        RECT 0.75 2.8 1.25 3.2 ;
      LAYER VIA12 ;
        RECT 0.87 2.87 1.13 3.13 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 2.75 3.65 3.25 ;
      LAYER MET2 ;
        RECT 3.3 2.75 3.7 3.25 ;
      LAYER VIA12 ;
        RECT 3.37 2.87 3.63 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 2.25 4.45 2.5 ;
        RECT 3.95 2.2 4.45 2.5 ;
        RECT 4.05 2.15 4.3 2.55 ;
        RECT 3.95 2.2 4.2 5.2 ;
        RECT 2.95 0.95 3.2 2.5 ;
      LAYER MET2 ;
        RECT 4 2.1 4.4 2.6 ;
      LAYER VIA12 ;
        RECT 4.07 2.22 4.33 2.48 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.1 3.75 3.35 5.2 ;
      RECT 1.4 3.75 1.65 5.2 ;
      RECT 1.4 3.75 3.35 4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi31_1

MACRO gf180mcu_osu_sc_gp9t3v3__buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_1 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 1.4 3.5 1.75 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 1.4 0 1.75 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.85 1.55 3.15 ;
      LAYER MET2 ;
        RECT 1.05 2.85 1.55 3.15 ;
        RECT 1.1 2.8 1.5 3.2 ;
      LAYER VIA12 ;
        RECT 1.17 2.87 1.43 3.13 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 3.5 2.75 3.8 ;
        RECT 2.45 1.5 2.7 3.8 ;
        RECT 2.35 3.5 2.6 5.2 ;
        RECT 2.35 0.95 2.6 1.8 ;
      LAYER MET2 ;
        RECT 2.25 3.45 2.75 3.85 ;
      LAYER VIA12 ;
        RECT 2.37 3.52 2.63 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.15 2.2 2.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_1

MACRO gf180mcu_osu_sc_gp9t3v3__buf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_16 0 0 ;
  SIZE 15.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15.8 6.15 ;
        RECT 15 3.5 15.25 6.15 ;
        RECT 13.3 3.5 13.55 6.15 ;
        RECT 11.6 3.5 11.85 6.15 ;
        RECT 9.9 3.5 10.15 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.05 3.5 14.55 3.8 ;
        RECT 14.15 0.95 14.4 5.2 ;
        RECT 2.25 2.95 14.4 3.25 ;
        RECT 2.25 2.05 14.4 2.35 ;
        RECT 12.45 0.95 12.7 5.2 ;
        RECT 10.75 0.95 11 5.2 ;
        RECT 9.05 0.95 9.3 5.2 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 14.05 3.45 14.55 3.85 ;
      LAYER VIA12 ;
        RECT 14.17 3.52 14.43 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_16

MACRO gf180mcu_osu_sc_gp9t3v3__buf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_2 0 0 ;
  SIZE 3.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.9 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 3.5 2.65 3.8 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 2.15 3.45 2.65 3.85 ;
      LAYER VIA12 ;
        RECT 2.27 3.52 2.53 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_2

MACRO gf180mcu_osu_sc_gp9t3v3__buf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_4 0 0 ;
  SIZE 5.65 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.65 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.65 0.6 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.85 3.5 4.35 3.8 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 2.95 4.2 3.25 ;
        RECT 2.25 2.05 4.2 2.35 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 3.85 3.45 4.35 3.85 ;
      LAYER VIA12 ;
        RECT 3.97 3.52 4.23 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_4

MACRO gf180mcu_osu_sc_gp9t3v3__buf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_8 0 0 ;
  SIZE 9.05 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 9.05 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.05 0.6 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 3.5 7.75 3.8 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 2.25 2.95 7.6 3.25 ;
        RECT 2.25 2.05 7.6 2.35 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 7.25 3.45 7.75 3.85 ;
      LAYER VIA12 ;
        RECT 7.37 3.52 7.63 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_8

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_1 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 1.4 3.5 1.75 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 1.4 0 1.75 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.85 1.55 3.15 ;
      LAYER MET2 ;
        RECT 1.05 2.85 1.55 3.15 ;
        RECT 1.1 2.8 1.5 3.2 ;
      LAYER VIA12 ;
        RECT 1.17 2.87 1.43 3.13 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 1.5 2.75 1.8 ;
        RECT 2.35 0.95 2.6 1.8 ;
        RECT 2.25 3.5 2.75 3.8 ;
        RECT 2.35 3.5 2.6 5.2 ;
      LAYER MET2 ;
        RECT 2.25 3.45 2.75 3.85 ;
        RECT 2.25 1.45 2.75 1.85 ;
        RECT 2.35 1.45 2.65 3.85 ;
      LAYER VIA12 ;
        RECT 2.37 3.52 2.63 3.78 ;
        RECT 2.37 1.52 2.63 1.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.15 2.2 2.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_1

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_16 0 0 ;
  SIZE 15.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15.8 6.15 ;
        RECT 15 3.5 15.25 6.15 ;
        RECT 13.3 3.5 13.55 6.15 ;
        RECT 11.6 3.5 11.85 6.15 ;
        RECT 9.9 3.5 10.15 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.05 3.5 14.55 3.8 ;
        RECT 14.15 0.95 14.4 5.2 ;
        RECT 2.25 2.95 14.4 3.25 ;
        RECT 2.25 2.05 14.4 2.35 ;
        RECT 12.45 0.95 12.7 5.2 ;
        RECT 10.75 0.95 11 5.2 ;
        RECT 9.05 0.95 9.3 5.2 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 14.05 3.45 14.55 3.85 ;
      LAYER VIA12 ;
        RECT 14.17 3.52 14.43 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_16

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_2 0 0 ;
  SIZE 3.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.9 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 3.5 2.65 3.8 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 2.15 3.45 2.65 3.85 ;
      LAYER VIA12 ;
        RECT 2.27 3.52 2.53 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_2

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_4 0 0 ;
  SIZE 5.65 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.65 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.65 0.6 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.85 3.5 4.35 3.8 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 2.95 4.2 3.25 ;
        RECT 2.25 2.05 4.2 2.35 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 3.85 3.45 4.35 3.85 ;
      LAYER VIA12 ;
        RECT 3.97 3.52 4.23 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_4

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_8 0 0 ;
  SIZE 9.05 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 9.05 6.15 ;
        RECT 8.2 3.5 8.45 6.15 ;
        RECT 6.5 3.5 6.75 6.15 ;
        RECT 4.8 3.5 5.05 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.05 0.6 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.2 1.55 2.5 ;
      LAYER MET2 ;
        RECT 1.05 2.2 1.55 2.5 ;
        RECT 1.1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.17 2.22 1.43 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.25 3.5 7.75 3.8 ;
        RECT 7.35 0.95 7.6 5.2 ;
        RECT 2.25 2.95 7.6 3.25 ;
        RECT 2.25 2.05 7.6 2.35 ;
        RECT 5.65 0.95 5.9 5.2 ;
        RECT 3.95 0.95 4.2 5.2 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 7.25 3.45 7.75 3.85 ;
      LAYER VIA12 ;
        RECT 7.37 3.52 7.63 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.95 2 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_8

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_1 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 0.55 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_1

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_16 0 0 ;
  SIZE 15 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15 6.15 ;
        RECT 14.15 3.5 14.4 6.15 ;
        RECT 12.45 3.5 12.7 6.15 ;
        RECT 10.75 3.5 11 6.15 ;
        RECT 9.05 3.5 9.3 6.15 ;
        RECT 7.35 3.5 7.6 6.15 ;
        RECT 5.65 3.5 5.9 6.15 ;
        RECT 3.95 3.5 4.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15 0.6 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 12.45 0 12.7 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 9.05 0 9.3 1.8 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.3 3.5 13.85 3.8 ;
        RECT 13.3 0.95 13.55 5.2 ;
        RECT 1.4 3 13.55 3.25 ;
        RECT 1.4 2.05 13.55 2.3 ;
        RECT 11.6 0.95 11.85 5.2 ;
        RECT 9.9 0.95 10.15 5.2 ;
        RECT 8.2 0.95 8.45 5.2 ;
        RECT 6.5 0.95 6.75 5.2 ;
        RECT 4.8 0.95 5.05 5.2 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 13.35 3.5 13.85 3.8 ;
        RECT 13.4 3.45 13.8 3.85 ;
      LAYER VIA12 ;
        RECT 13.47 3.52 13.73 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_16

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_2 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 2.3 3.5 2.55 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 2.2 1.15 2.5 ;
      LAYER MET2 ;
        RECT 0.65 2.15 1.15 2.55 ;
      LAYER VIA12 ;
        RECT 0.77 2.22 1.03 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 3.5 2.05 3.8 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.55 3.5 2.05 3.8 ;
        RECT 1.6 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.67 3.52 1.93 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_2

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_4 0 0 ;
  SIZE 4.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.8 6.15 ;
        RECT 4 3.5 4.25 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 3.5 3.75 3.8 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 3 3.35 3.25 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 3.25 3.5 3.75 3.8 ;
        RECT 3.3 3.45 3.7 3.85 ;
      LAYER VIA12 ;
        RECT 3.37 3.52 3.63 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_4

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_8 0 0 ;
  SIZE 8.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.2 6.15 ;
        RECT 7.4 3.5 7.65 6.15 ;
        RECT 5.65 3.5 5.9 6.15 ;
        RECT 3.95 3.5 4.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.2 0.6 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.5 3.5 7.15 3.8 ;
        RECT 6.5 0.95 6.75 5.2 ;
        RECT 1.4 3 6.75 3.25 ;
        RECT 1.4 2.05 6.75 2.3 ;
        RECT 4.8 0.95 5.05 5.2 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 6.65 3.5 7.15 3.8 ;
        RECT 6.7 3.45 7.1 3.85 ;
      LAYER VIA12 ;
        RECT 6.77 3.52 7.03 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_8

MACRO gf180mcu_osu_sc_gp9t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dff_1 0 0 ;
  SIZE 14.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 14.5 6.15 ;
        RECT 12.85 4.05 13.1 6.15 ;
        RECT 10.4 3.5 10.65 6.15 ;
        RECT 8.6 4.75 8.85 6.15 ;
        RECT 5 4.1 5.25 6.15 ;
        RECT 1.4 4.75 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.5 0.6 ;
        RECT 12.85 0 13.1 1.6 ;
        RECT 10.4 0 10.65 1.4 ;
        RECT 8.6 0 8.85 1.5 ;
        RECT 5 0 5.25 1.4 ;
        RECT 1.4 0 1.65 1.5 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 2.5 3 9.4 3.25 ;
        RECT 2.5 3 8.95 3.3 ;
        RECT 5.95 1.95 6.45 2.25 ;
        RECT 6.05 1.95 6.35 3.3 ;
        RECT 3.8 2 4.3 2.3 ;
        RECT 3.9 2 4.2 3.3 ;
      LAYER MET2 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 9.05 2.8 9.45 3.2 ;
      LAYER VIA12 ;
        RECT 9.12 2.87 9.38 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 2.85 2.25 3.15 ;
      LAYER MET2 ;
        RECT 1.7 2.85 2.3 3.15 ;
        RECT 1.75 2.8 2.25 3.2 ;
      LAYER VIA12 ;
        RECT 1.87 2.87 2.13 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.7 4.15 14.25 4.5 ;
        RECT 13.7 4.1 14.2 4.5 ;
        RECT 13.7 0.95 13.95 5.2 ;
      LAYER MET2 ;
        RECT 13.75 4.15 14.25 4.45 ;
        RECT 13.8 4.1 14.2 4.5 ;
      LAYER VIA12 ;
        RECT 13.87 4.17 14.13 4.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12 3.5 13.45 3.8 ;
        RECT 13.05 1.85 13.35 3.8 ;
        RECT 12 1.85 13.35 2.1 ;
        RECT 12 3.5 12.25 5.2 ;
        RECT 12 0.95 12.25 2.1 ;
      LAYER MET2 ;
        RECT 12.95 3.5 13.45 3.8 ;
        RECT 13 3.45 13.4 3.85 ;
      LAYER VIA12 ;
        RECT 13.07 3.52 13.33 3.78 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 8.1 4.15 8.5 4.55 ;
      RECT 8.05 4.2 11.45 4.5 ;
      RECT 11.15 2.55 11.45 4.5 ;
      RECT 8.15 2.15 8.45 4.55 ;
      RECT 12.2 2.5 12.6 2.9 ;
      RECT 11.15 2.55 12.65 2.85 ;
      RECT 8.1 2.15 8.5 2.55 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 6.4 0.9 6.7 4.6 ;
      RECT 6.35 4.15 6.75 4.55 ;
      RECT 10.55 1.6 10.95 2 ;
      RECT 10.2 1.65 11 1.95 ;
      RECT 6.35 1.3 6.75 1.7 ;
      RECT 6.4 0.9 6.75 1.7 ;
      RECT 6.3 1.35 6.75 1.65 ;
      RECT 10.2 1.6 10.95 1.95 ;
      RECT 10.2 0.9 10.5 1.95 ;
      RECT 6.4 0.9 10.5 1.2 ;
      RECT 2.8 4.9 7.55 5.2 ;
      RECT 7.25 1.5 7.55 5.2 ;
      RECT 2.8 1.95 3.1 5.2 ;
      RECT 2.75 1.95 3.2 2.35 ;
      RECT 2.7 2 3.2 2.3 ;
      RECT 9.4 1.5 9.8 1.9 ;
      RECT 7.2 1.5 7.6 1.9 ;
      RECT 7.15 1.55 9.9 1.85 ;
      RECT 4.65 1.95 5.05 2.35 ;
      RECT 0.45 1.95 0.85 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 0.4 2 0.9 2.3 ;
      RECT 4.7 1.05 5 2.35 ;
      RECT 0.5 1.05 0.8 2.35 ;
      RECT 0.5 1.05 5 1.35 ;
    LAYER VIA12 ;
      RECT 12.27 2.57 12.53 2.83 ;
      RECT 10.62 1.67 10.88 1.93 ;
      RECT 9.47 1.57 9.73 1.83 ;
      RECT 8.17 2.22 8.43 2.48 ;
      RECT 8.17 4.22 8.43 4.48 ;
      RECT 7.27 1.57 7.53 1.83 ;
      RECT 6.42 1.37 6.68 1.63 ;
      RECT 6.42 4.22 6.68 4.48 ;
      RECT 4.72 2.02 4.98 2.28 ;
      RECT 2.82 2.02 3.08 2.28 ;
      RECT 0.52 2.02 0.78 2.28 ;
    LAYER MET1 ;
      RECT 11.25 0.95 11.5 5.2 ;
      RECT 11.25 2.55 12.65 2.85 ;
      RECT 10.6 1.65 10.9 2.95 ;
      RECT 10.5 1.65 11 1.95 ;
      RECT 9.45 3.5 9.7 5.2 ;
      RECT 9.45 3.5 10 3.75 ;
      RECT 9.75 2.2 10 3.75 ;
      RECT 9.45 1.45 9.75 2.5 ;
      RECT 9.45 0.95 9.7 2.5 ;
      RECT 8.05 4.2 8.55 4.5 ;
      RECT 8.15 4.1 8.45 4.5 ;
      RECT 6.95 1.9 7.25 2.4 ;
      RECT 6.9 2 7.55 2.3 ;
      RECT 7.25 1.45 7.55 2.3 ;
      RECT 6.3 1.4 6.95 1.65 ;
      RECT 6.4 0.95 6.95 1.65 ;
      RECT 6.4 4.2 6.95 5.2 ;
      RECT 6.4 4.1 6.7 5.2 ;
      RECT 4.7 2 5 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 3.3 4.2 3.85 5.2 ;
      RECT 1.05 4.2 3.85 4.5 ;
      RECT 1.05 1.8 1.35 4.5 ;
      RECT 1.05 3 1.45 3.3 ;
      RECT 1.05 1.8 2.25 2.05 ;
      RECT 2 1.4 2.25 2.05 ;
      RECT 2 1.4 3.85 1.65 ;
      RECT 3.3 0.95 3.85 1.65 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.5 1.9 0.8 2.35 ;
      RECT 0.4 2 0.8 2.3 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 2.7 2 3.2 2.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dff_1

MACRO gf180mcu_osu_sc_gp9t3v3__dffn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffn_1 0 0 ;
  SIZE 14.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 14.5 6.15 ;
        RECT 12.85 4.05 13.1 6.15 ;
        RECT 10.4 3.5 10.65 6.15 ;
        RECT 8.6 4.75 8.85 6.15 ;
        RECT 5 4.1 5.25 6.15 ;
        RECT 1.4 4.75 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.5 0.6 ;
        RECT 12.85 0 13.1 1.6 ;
        RECT 10.4 0 10.65 1.4 ;
        RECT 8.6 0 8.85 1.5 ;
        RECT 5 0 5.25 1.4 ;
        RECT 1.4 0 1.65 1.5 ;
    END
  END VSS
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 2.5 3 9.4 3.25 ;
        RECT 2.5 3 8.95 3.3 ;
        RECT 5.95 1.95 6.45 2.25 ;
        RECT 6.05 1.95 6.35 3.3 ;
        RECT 3.8 2 4.3 2.3 ;
        RECT 3.9 2 4.2 3.3 ;
      LAYER MET2 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 9.05 2.8 9.45 3.2 ;
      LAYER VIA12 ;
        RECT 9.12 2.87 9.38 3.13 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 2.85 2.25 3.15 ;
      LAYER MET2 ;
        RECT 1.7 2.85 2.3 3.15 ;
        RECT 1.75 2.8 2.25 3.2 ;
      LAYER VIA12 ;
        RECT 1.87 2.87 2.13 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.7 4.15 14.25 4.5 ;
        RECT 13.7 4.1 14.2 4.5 ;
        RECT 13.7 0.95 13.95 5.2 ;
      LAYER MET2 ;
        RECT 13.75 4.15 14.25 4.45 ;
        RECT 13.8 4.1 14.2 4.5 ;
      LAYER VIA12 ;
        RECT 13.87 4.17 14.13 4.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12 3.5 13.45 3.8 ;
        RECT 13.05 1.85 13.35 3.8 ;
        RECT 12 1.85 13.35 2.1 ;
        RECT 12 3.5 12.25 5.2 ;
        RECT 12 0.95 12.25 2.1 ;
      LAYER MET2 ;
        RECT 12.95 3.5 13.45 3.8 ;
        RECT 13 3.45 13.4 3.85 ;
      LAYER VIA12 ;
        RECT 13.07 3.52 13.33 3.78 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 8.1 4.15 8.5 4.55 ;
      RECT 8.05 4.2 11.45 4.5 ;
      RECT 11.15 2.55 11.45 4.5 ;
      RECT 8.15 2.15 8.45 4.55 ;
      RECT 12.2 2.5 12.6 2.9 ;
      RECT 11.15 2.55 12.65 2.85 ;
      RECT 8.1 2.15 8.5 2.55 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 6.4 0.9 6.7 4.6 ;
      RECT 6.35 4.15 6.75 4.55 ;
      RECT 10.55 1.6 10.95 2 ;
      RECT 10.2 1.65 11 1.95 ;
      RECT 6.35 1.3 6.75 1.7 ;
      RECT 6.4 0.9 6.75 1.7 ;
      RECT 6.3 1.35 6.75 1.65 ;
      RECT 10.2 1.6 10.95 1.95 ;
      RECT 10.2 0.9 10.5 1.95 ;
      RECT 6.4 0.9 10.5 1.2 ;
      RECT 2.8 4.9 7.55 5.2 ;
      RECT 7.25 1.5 7.55 5.2 ;
      RECT 2.8 1.95 3.1 5.2 ;
      RECT 2.75 1.95 3.2 2.35 ;
      RECT 2.7 2 3.2 2.3 ;
      RECT 9.4 1.5 9.8 1.9 ;
      RECT 7.2 1.5 7.6 1.9 ;
      RECT 7.15 1.55 9.9 1.85 ;
      RECT 4.65 1.95 5.05 2.35 ;
      RECT 0.45 1.95 0.85 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 0.4 2 0.9 2.3 ;
      RECT 4.7 1.05 5 2.35 ;
      RECT 0.5 1.05 0.8 2.35 ;
      RECT 0.5 1.05 5 1.35 ;
    LAYER VIA12 ;
      RECT 12.27 2.57 12.53 2.83 ;
      RECT 10.62 1.67 10.88 1.93 ;
      RECT 9.47 1.57 9.73 1.83 ;
      RECT 8.17 2.22 8.43 2.48 ;
      RECT 8.17 4.22 8.43 4.48 ;
      RECT 7.27 1.57 7.53 1.83 ;
      RECT 6.42 1.37 6.68 1.63 ;
      RECT 6.42 4.22 6.68 4.48 ;
      RECT 4.72 2.02 4.98 2.28 ;
      RECT 2.82 2.02 3.08 2.28 ;
      RECT 0.52 2.02 0.78 2.28 ;
    LAYER MET1 ;
      RECT 11.25 0.95 11.5 5.2 ;
      RECT 11.25 2.55 12.65 2.85 ;
      RECT 10.6 1.65 10.9 2.95 ;
      RECT 10.5 1.65 11 1.95 ;
      RECT 9.45 3.5 9.7 5.2 ;
      RECT 9.45 3.5 10 3.75 ;
      RECT 9.75 2.2 10 3.75 ;
      RECT 9.45 1.45 9.75 2.5 ;
      RECT 9.45 0.95 9.7 2.5 ;
      RECT 8.05 4.2 8.55 4.5 ;
      RECT 8.15 4.1 8.45 4.5 ;
      RECT 6.95 1.9 7.25 2.4 ;
      RECT 6.9 2 7.55 2.3 ;
      RECT 7.25 1.45 7.55 2.3 ;
      RECT 6.3 1.4 6.95 1.65 ;
      RECT 6.4 0.95 6.95 1.65 ;
      RECT 6.4 4.2 6.95 5.2 ;
      RECT 6.4 4.1 6.7 5.2 ;
      RECT 4.7 2 5 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 3.3 4.2 3.85 5.2 ;
      RECT 1.05 4.2 3.85 4.5 ;
      RECT 1.05 1.8 1.35 4.5 ;
      RECT 1.05 3 1.45 3.3 ;
      RECT 1.05 1.8 2.25 2.05 ;
      RECT 2 1.4 2.25 2.05 ;
      RECT 2 1.4 3.85 1.65 ;
      RECT 3.3 0.95 3.85 1.65 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.5 1.9 0.8 2.35 ;
      RECT 0.4 2 0.8 2.3 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 2.7 2 3.2 2.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffn_1

MACRO gf180mcu_osu_sc_gp9t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffsr_1 0 0 ;
  SIZE 20.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 20.5 6.15 ;
        RECT 18.8 4.05 19.05 6.15 ;
        RECT 15.5 4.25 15.75 6.15 ;
        RECT 12.9 4.75 13.15 6.15 ;
        RECT 9.3 4.1 9.55 6.15 ;
        RECT 5.7 4.75 5.95 6.15 ;
        RECT 3.85 4.25 4.1 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 20.5 0.6 ;
        RECT 18.8 0 19.05 1.6 ;
        RECT 17.05 0 17.3 1.4 ;
        RECT 14.8 0 15.05 1.8 ;
        RECT 12.9 0 13.15 1.7 ;
        RECT 9.3 0 9.55 1.4 ;
        RECT 5.7 0 5.95 1.5 ;
        RECT 4.55 0 4.8 1.45 ;
        RECT 2.3 0 2.55 1.4 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 13.3 2.85 13.8 3.15 ;
        RECT 6.8 3 13.7 3.3 ;
        RECT 10.25 2.2 10.75 2.45 ;
        RECT 10.35 2.2 10.65 3.3 ;
        RECT 8.1 2.15 8.6 2.45 ;
        RECT 8.2 2.15 8.5 3.3 ;
      LAYER MET2 ;
        RECT 13.3 2.85 13.8 3.15 ;
        RECT 13.35 2.8 13.75 3.2 ;
      LAYER VIA12 ;
        RECT 13.42 2.87 13.68 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.05 2.85 6.55 3.15 ;
      LAYER MET2 ;
        RECT 6 2.85 6.6 3.15 ;
        RECT 6.05 2.8 6.55 3.2 ;
      LAYER VIA12 ;
        RECT 6.17 2.87 6.43 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 19.65 0.95 19.9 5.2 ;
        RECT 19.6 4.05 19.9 4.55 ;
      LAYER MET2 ;
        RECT 19.5 4.15 20 4.45 ;
        RECT 19.55 4.1 19.95 4.5 ;
      LAYER VIA12 ;
        RECT 19.62 4.17 19.88 4.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 17.95 3.5 19.4 3.8 ;
        RECT 19 3.45 19.3 3.8 ;
        RECT 19.05 1.85 19.3 3.8 ;
        RECT 17.95 1.85 19.3 2.1 ;
        RECT 17.95 3.5 18.2 5.2 ;
        RECT 17.95 0.95 18.2 2.1 ;
      LAYER MET2 ;
        RECT 18.9 3.5 19.4 3.8 ;
        RECT 18.95 3.45 19.35 3.85 ;
      LAYER VIA12 ;
        RECT 19.02 3.52 19.28 3.78 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.8 2.75 1.1 3.25 ;
      LAYER MET2 ;
        RECT 0.7 2.85 1.2 3.15 ;
        RECT 0.75 2.8 1.15 3.2 ;
      LAYER VIA12 ;
        RECT 0.82 2.87 1.08 3.13 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.9 2.85 16.4 3.15 ;
        RECT 3.4 3 3.9 3.3 ;
      LAYER MET2 ;
        RECT 15.9 2.8 16.4 3.2 ;
        RECT 3.5 4.95 16.3 5.25 ;
        RECT 16 2.8 16.3 5.25 ;
        RECT 3.4 2.95 3.9 3.35 ;
        RECT 3.5 2.95 3.8 5.25 ;
      LAYER VIA12 ;
        RECT 3.52 3.02 3.78 3.28 ;
        RECT 16.02 2.87 16.28 3.13 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 18.15 2.5 18.55 2.9 ;
      RECT 18 2.55 18.6 2.85 ;
      RECT 16.6 2.05 16.9 2.55 ;
      RECT 2.65 2.15 3.15 2.55 ;
      RECT 1.35 2.15 1.75 2.55 ;
      RECT 16.55 2.05 16.95 2.5 ;
      RECT 1.3 2.2 3.15 2.5 ;
      RECT 2.75 0.9 3.05 2.55 ;
      RECT 16.55 0.9 16.85 2.5 ;
      RECT 2.75 0.9 16.85 1.2 ;
      RECT 10.7 1.5 11 4.05 ;
      RECT 10.65 3.6 11.05 4 ;
      RECT 14.6 2 15.1 2.4 ;
      RECT 14.6 1.55 15 2.4 ;
      RECT 10.65 1.5 11.05 1.9 ;
      RECT 10.6 1.55 15 1.85 ;
      RECT 12.4 4.15 12.8 4.55 ;
      RECT 12.35 4.2 14.5 4.5 ;
      RECT 14.2 2.85 14.5 4.5 ;
      RECT 12.45 2.4 12.75 4.55 ;
      RECT 14.2 2.85 15.05 3.2 ;
      RECT 14.55 2.8 15.05 3.2 ;
      RECT 12.4 2.4 12.8 2.8 ;
      RECT 12.35 2.45 12.85 2.75 ;
      RECT 7.1 4.35 11.7 4.65 ;
      RECT 11.4 2.15 11.7 4.65 ;
      RECT 7.1 2.1 7.4 4.65 ;
      RECT 11.35 2.2 11.75 2.6 ;
      RECT 7.05 2.1 7.5 2.5 ;
      RECT 7 2.15 7.5 2.45 ;
      RECT 9 1.5 9.3 2.4 ;
      RECT 8.95 1.95 9.35 2.35 ;
      RECT 8.95 2 9.4 2.3 ;
      RECT 4.65 1.85 5.15 2.25 ;
      RECT 4.65 1.9 6.6 2.2 ;
      RECT 6.3 1.5 6.6 2.2 ;
      RECT 8.95 1.5 9.3 2.35 ;
      RECT 6.3 1.5 9.3 1.8 ;
      RECT 4.4 2.95 4.9 3.35 ;
    LAYER VIA12 ;
      RECT 18.22 2.57 18.48 2.83 ;
      RECT 16.62 2.17 16.88 2.43 ;
      RECT 14.72 2.07 14.98 2.33 ;
      RECT 14.67 2.87 14.93 3.13 ;
      RECT 12.47 2.47 12.73 2.73 ;
      RECT 12.47 4.22 12.73 4.48 ;
      RECT 11.42 2.27 11.68 2.53 ;
      RECT 10.72 1.57 10.98 1.83 ;
      RECT 10.72 3.67 10.98 3.93 ;
      RECT 9.02 2.02 9.28 2.28 ;
      RECT 7.12 2.17 7.38 2.43 ;
      RECT 4.77 1.92 5.03 2.18 ;
      RECT 4.52 3.02 4.78 3.28 ;
      RECT 2.77 2.22 3.03 2.48 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 17.2 3.85 17.45 5.2 ;
      RECT 17.25 1.65 17.5 4.1 ;
      RECT 14.55 2.85 15.65 3.15 ;
      RECT 15.35 1.65 15.65 3.15 ;
      RECT 17.25 2.55 18.6 2.85 ;
      RECT 15.35 1.65 17.5 1.9 ;
      RECT 16.2 0.95 16.45 1.9 ;
      RECT 16.35 3.75 16.6 5.2 ;
      RECT 14.65 3.75 14.9 5.2 ;
      RECT 14.65 3.75 16.6 4 ;
      RECT 13.75 3.6 14 5.2 ;
      RECT 13.75 3.6 14.3 3.85 ;
      RECT 14.05 2.2 14.3 3.85 ;
      RECT 11.4 1.95 11.7 2.7 ;
      RECT 13.75 2.2 14.3 2.5 ;
      RECT 11.4 1.95 14 2.2 ;
      RECT 13.75 0.95 14 2.5 ;
      RECT 12.35 4.2 12.85 4.5 ;
      RECT 12.45 4.1 12.75 4.5 ;
      RECT 10.7 0.95 11 1.95 ;
      RECT 10.7 0.95 11.25 1.65 ;
      RECT 10.7 3.7 11.25 5.2 ;
      RECT 10.7 3.55 11 5.2 ;
      RECT 9 2 9.3 2.35 ;
      RECT 8.9 2 9.4 2.3 ;
      RECT 7.6 4.2 8.15 5.2 ;
      RECT 5.4 4.2 8.15 4.5 ;
      RECT 5.4 2.2 5.7 4.5 ;
      RECT 4.4 3 5.7 3.3 ;
      RECT 5.4 2.2 6.55 2.5 ;
      RECT 6.25 1.4 6.55 2.5 ;
      RECT 6.25 1.4 8.15 1.65 ;
      RECT 7.6 0.95 8.15 1.65 ;
      RECT 2.15 1.65 2.4 5.2 ;
      RECT 3.85 1.9 5.15 2.2 ;
      RECT 3.15 1.6 4.1 1.9 ;
      RECT 2.15 1.65 4.1 1.9 ;
      RECT 3.15 0.95 3.4 1.9 ;
      RECT 4.7 3.75 4.95 5.2 ;
      RECT 3 3.75 3.25 5.2 ;
      RECT 3 3.75 4.95 4 ;
      RECT 1.4 0.95 1.65 5.2 ;
      RECT 1.4 1.9 1.7 2.55 ;
      RECT 1.4 2.2 1.8 2.5 ;
      RECT 16.5 2.15 17 2.45 ;
      RECT 14.6 2.05 15.1 2.35 ;
      RECT 12.35 2.45 12.85 2.75 ;
      RECT 7 2.15 7.5 2.45 ;
      RECT 2.65 2.2 3.15 2.5 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffsr_1

MACRO gf180mcu_osu_sc_gp9t3v3__dlat_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlat_1 0 0 ;
  SIZE 9.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 9.5 6.15 ;
        RECT 7.8 4.2 8.05 6.15 ;
        RECT 5.35 3.75 5.6 6.15 ;
        RECT 1.45 4.3 1.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.5 0.6 ;
        RECT 7.8 0 8.05 1.45 ;
        RECT 5.2 0 5.6 1.45 ;
        RECT 1.45 0 1.85 1.5 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 5.7 3 6.2 3.3 ;
        RECT 3.4 2.85 3.9 3.3 ;
      LAYER MET2 ;
        RECT 5.7 2.95 6.2 3.35 ;
        RECT 3.5 3 6.2 3.3 ;
        RECT 3.4 2.85 3.9 3.15 ;
        RECT 3.45 2.8 3.85 3.2 ;
      LAYER VIA12 ;
        RECT 3.52 2.87 3.78 3.13 ;
        RECT 5.82 3.02 6.08 3.28 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.65 2.85 9.15 3.15 ;
        RECT 8.65 2.8 9.05 3.2 ;
        RECT 8.65 0.95 8.9 5.2 ;
      LAYER MET2 ;
        RECT 8.65 2.85 9.15 3.15 ;
        RECT 8.7 2.8 9.1 3.2 ;
      LAYER VIA12 ;
        RECT 8.77 2.87 9.03 3.13 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 7.2 2.3 7.7 2.7 ;
      RECT 5.05 2.3 5.45 2.7 ;
      RECT 4.6 2.35 7.7 2.65 ;
      RECT 0.35 2.15 0.85 2.55 ;
      RECT 0.35 2.2 4.9 2.5 ;
      RECT 0.35 2.3 5.45 2.5 ;
    LAYER VIA12 ;
      RECT 7.32 2.37 7.58 2.63 ;
      RECT 5.12 2.37 5.38 2.63 ;
      RECT 0.47 2.22 0.73 2.48 ;
    LAYER MET1 ;
      RECT 6.95 3.35 7.2 5.2 ;
      RECT 6.95 3.35 8.3 3.6 ;
      RECT 8 1.85 8.3 3.6 ;
      RECT 6.95 1.85 8.3 2.1 ;
      RECT 6.95 0.95 7.2 2.1 ;
      RECT 6.2 3.65 6.45 5.2 ;
      RECT 6.45 2 6.7 3.9 ;
      RECT 2.6 3 3.1 3.3 ;
      RECT 2.7 2.3 3 3.3 ;
      RECT 4.15 2.45 4.65 2.75 ;
      RECT 2.7 2.3 4.5 2.6 ;
      RECT 2.7 2.35 4.55 2.6 ;
      RECT 4.2 1.7 4.5 2.75 ;
      RECT 6.2 0.95 6.45 2.25 ;
      RECT 4.2 1.7 6.45 1.95 ;
      RECT 3.15 3.8 3.4 5.2 ;
      RECT 1.15 3.8 3.4 4.05 ;
      RECT 1.15 1.9 1.4 4.05 ;
      RECT 1.1 3 1.55 3.3 ;
      RECT 1.15 1.9 2.4 2.15 ;
      RECT 2.15 1.2 2.4 2.15 ;
      RECT 3.15 0.95 3.4 1.55 ;
      RECT 2.15 1.2 3.4 1.45 ;
      RECT 0.6 0.95 0.85 5.2 ;
      RECT 0.5 2.15 0.85 2.55 ;
      RECT 0.35 2.2 0.85 2.5 ;
      RECT 0.45 2.15 0.85 2.5 ;
      RECT 7.2 2.35 7.7 2.65 ;
      RECT 5 2.35 5.5 2.65 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlat_1

MACRO gf180mcu_osu_sc_gp9t3v3__dlatn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dlatn_1 0 0 ;
  SIZE 9.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 9.5 6.15 ;
        RECT 7.8 4.2 8.05 6.15 ;
        RECT 5.35 3.75 5.6 6.15 ;
        RECT 1.45 4.3 1.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 9.5 0.6 ;
        RECT 7.8 0 8.05 1.45 ;
        RECT 5.2 0 5.6 1.45 ;
        RECT 1.45 0 1.85 1.5 ;
    END
  END VSS
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 5.7 3 6.2 3.3 ;
        RECT 3.4 2.85 3.9 3.3 ;
      LAYER MET2 ;
        RECT 5.7 2.95 6.2 3.35 ;
        RECT 3.5 3 6.2 3.3 ;
        RECT 3.4 2.85 3.9 3.15 ;
        RECT 3.45 2.8 3.85 3.2 ;
      LAYER VIA12 ;
        RECT 3.52 2.87 3.78 3.13 ;
        RECT 5.82 3.02 6.08 3.28 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.65 2.85 9.15 3.15 ;
        RECT 8.65 2.8 9.05 3.2 ;
        RECT 8.65 0.95 8.9 5.2 ;
      LAYER MET2 ;
        RECT 8.65 2.85 9.15 3.15 ;
        RECT 8.7 2.8 9.1 3.2 ;
      LAYER VIA12 ;
        RECT 8.77 2.87 9.03 3.13 ;
    END
  END Q
  OBS
    LAYER MET2 ;
      RECT 7.2 2.3 7.7 2.7 ;
      RECT 5.05 2.3 5.45 2.7 ;
      RECT 4.6 2.35 7.7 2.65 ;
      RECT 0.35 2.15 0.85 2.55 ;
      RECT 0.35 2.2 4.9 2.5 ;
      RECT 0.35 2.3 5.45 2.5 ;
    LAYER VIA12 ;
      RECT 7.32 2.37 7.58 2.63 ;
      RECT 5.12 2.37 5.38 2.63 ;
      RECT 0.47 2.22 0.73 2.48 ;
    LAYER MET1 ;
      RECT 6.95 3.35 7.2 5.2 ;
      RECT 6.95 3.35 8.3 3.6 ;
      RECT 8 1.85 8.3 3.6 ;
      RECT 6.95 1.85 8.3 2.1 ;
      RECT 6.95 0.95 7.2 2.1 ;
      RECT 6.2 3.65 6.45 5.2 ;
      RECT 6.45 2 6.7 3.9 ;
      RECT 2.6 3 3.1 3.3 ;
      RECT 2.7 2.3 3 3.3 ;
      RECT 4.15 2.45 4.65 2.75 ;
      RECT 2.7 2.3 4.5 2.6 ;
      RECT 2.7 2.35 4.55 2.6 ;
      RECT 4.2 1.7 4.5 2.75 ;
      RECT 6.2 0.95 6.45 2.25 ;
      RECT 4.2 1.7 6.45 1.95 ;
      RECT 3.15 3.8 3.4 5.2 ;
      RECT 1.15 3.8 3.4 4.05 ;
      RECT 1.15 1.9 1.4 4.05 ;
      RECT 1.1 3 1.55 3.3 ;
      RECT 1.15 1.9 2.4 2.15 ;
      RECT 2.15 1.2 2.4 2.15 ;
      RECT 3.15 0.95 3.4 1.55 ;
      RECT 2.15 1.2 3.4 1.45 ;
      RECT 0.6 0.95 0.85 5.2 ;
      RECT 0.5 2.15 0.85 2.55 ;
      RECT 0.35 2.2 0.85 2.5 ;
      RECT 0.45 2.15 0.85 2.5 ;
      RECT 7.2 2.35 7.7 2.65 ;
      RECT 5 2.35 5.5 2.65 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dlatn_1

MACRO gf180mcu_osu_sc_gp9t3v3__fill_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_1 0 0 ;
  SIZE 0.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 0.1 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.1 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__fill_1

MACRO gf180mcu_osu_sc_gp9t3v3__fill_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_16 0 0 ;
  SIZE 1.6 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 1.6 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 1.6 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__fill_16

MACRO gf180mcu_osu_sc_gp9t3v3__fill_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_2 0 0 ;
  SIZE 0.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 0.2 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.2 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__fill_2

MACRO gf180mcu_osu_sc_gp9t3v3__fill_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_4 0 0 ;
  SIZE 0.4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 0.4 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.4 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__fill_4

MACRO gf180mcu_osu_sc_gp9t3v3__fill_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__fill_8 0 0 ;
  SIZE 0.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 0.8 0.6 ;
    END
  END VSS
END gf180mcu_osu_sc_gp9t3v3__fill_8

MACRO gf180mcu_osu_sc_gp9t3v3__inv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_1 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 0.55 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_1

MACRO gf180mcu_osu_sc_gp9t3v3__inv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_16 0 0 ;
  SIZE 15 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15 6.15 ;
        RECT 14.15 3.5 14.4 6.15 ;
        RECT 12.45 3.5 12.7 6.15 ;
        RECT 10.75 3.5 11 6.15 ;
        RECT 9.05 3.5 9.3 6.15 ;
        RECT 7.35 3.5 7.6 6.15 ;
        RECT 5.65 3.5 5.9 6.15 ;
        RECT 3.95 3.5 4.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15 0.6 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 12.45 0 12.7 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 9.05 0 9.3 1.8 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.3 3.5 13.85 3.8 ;
        RECT 13.3 0.95 13.55 5.2 ;
        RECT 1.4 3 13.55 3.25 ;
        RECT 1.4 2.05 13.55 2.3 ;
        RECT 11.6 0.95 11.85 5.2 ;
        RECT 9.9 0.95 10.15 5.2 ;
        RECT 8.2 0.95 8.45 5.2 ;
        RECT 6.5 0.95 6.75 5.2 ;
        RECT 4.8 0.95 5.05 5.2 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 13.35 3.5 13.85 3.8 ;
        RECT 13.4 3.45 13.8 3.85 ;
      LAYER VIA12 ;
        RECT 13.47 3.52 13.73 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_16

MACRO gf180mcu_osu_sc_gp9t3v3__inv_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_2 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 2.3 3.5 2.55 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.65 2.2 1.15 2.5 ;
      LAYER MET2 ;
        RECT 0.65 2.15 1.15 2.55 ;
      LAYER VIA12 ;
        RECT 0.77 2.22 1.03 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 3.5 2.05 3.8 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.55 3.5 2.05 3.8 ;
        RECT 1.6 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.67 3.52 1.93 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_2

MACRO gf180mcu_osu_sc_gp9t3v3__inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_4 0 0 ;
  SIZE 4.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.8 6.15 ;
        RECT 4 3.5 4.25 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 3.5 3.75 3.8 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 3 3.35 3.25 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 3.25 3.5 3.75 3.8 ;
        RECT 3.3 3.45 3.7 3.85 ;
      LAYER VIA12 ;
        RECT 3.37 3.52 3.63 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_4

MACRO gf180mcu_osu_sc_gp9t3v3__inv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_8 0 0 ;
  SIZE 8.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.2 6.15 ;
        RECT 7.4 3.5 7.65 6.15 ;
        RECT 5.65 3.5 5.9 6.15 ;
        RECT 3.95 3.5 4.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.2 0.6 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.5 3.5 7.15 3.8 ;
        RECT 6.5 0.95 6.75 5.2 ;
        RECT 1.4 3 6.75 3.25 ;
        RECT 1.4 2.05 6.75 2.3 ;
        RECT 4.8 0.95 5.05 5.2 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 6.65 3.5 7.15 3.8 ;
        RECT 6.7 3.45 7.1 3.85 ;
      LAYER VIA12 ;
        RECT 6.77 3.52 7.03 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_8

MACRO gf180mcu_osu_sc_gp9t3v3__lshifdown
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__lshifdown 0 0 ;
  SIZE 4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 2.15 5.55 4 6.15 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 1.85 6.15 ;
        RECT 0.55 3.5 0.85 6.15 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4 0.6 ;
        RECT 2.25 0 2.55 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 0.55 2.15 1.05 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 2.2 3.5 2.5 ;
        RECT 3.15 0.95 3.45 5.2 ;
      LAYER MET2 ;
        RECT 3.05 2.15 3.55 2.55 ;
      LAYER VIA12 ;
        RECT 3.17 2.22 3.43 2.48 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.3 2.8 2.8 3.2 ;
      RECT 1.45 2.85 2.8 3.15 ;
      RECT 1.45 2.15 1.75 3.15 ;
      RECT 1.35 2.15 1.85 2.55 ;
    LAYER VIA12 ;
      RECT 2.42 2.87 2.68 3.13 ;
      RECT 1.47 2.22 1.73 2.48 ;
    LAYER MET1 ;
      RECT 1.45 0.95 1.75 5.2 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 2.3 2.85 2.8 3.15 ;
      RECT 2.25 3.5 2.55 5.2 ;
  END
END gf180mcu_osu_sc_gp9t3v3__lshifdown

MACRO gf180mcu_osu_sc_gp9t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__lshifup 0 0 ;
  SIZE 7.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 1.9 6.15 ;
        RECT 0.55 3.5 0.85 6.15 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.15 5.55 7.1 6.15 ;
        RECT 5.35 3.5 5.65 6.15 ;
        RECT 3.3 4.05 3.8 6.15 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 7.1 0.6 ;
        RECT 5.35 0 5.65 1.8 ;
        RECT 3.3 0 3.8 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.65 2.05 3.15 2.35 ;
        RECT 0.55 2.2 1.05 2.5 ;
      LAYER MET2 ;
        RECT 2.65 2.05 3.15 2.35 ;
        RECT 2.65 2 3.1 2.4 ;
        RECT 2.8 1.4 3.1 2.4 ;
        RECT 0.7 1.4 3.1 1.7 ;
        RECT 0.55 2.15 1.05 2.55 ;
        RECT 0.7 1.4 1 2.55 ;
      LAYER VIA12 ;
        RECT 0.67 2.22 0.93 2.48 ;
        RECT 2.77 2.07 3.03 2.33 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.2 2.2 6.6 2.5 ;
        RECT 6.25 0.95 6.55 5.2 ;
      LAYER MET2 ;
        RECT 6.15 2.15 6.65 2.55 ;
      LAYER VIA12 ;
        RECT 6.27 2.22 6.53 2.48 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.2 3.5 2.7 3.9 ;
      RECT 2.2 3.5 4.45 3.85 ;
      RECT 4.15 2.8 4.45 3.85 ;
      RECT 5.4 2.8 5.9 3.2 ;
      RECT 4.1 2.8 4.5 3.2 ;
      RECT 4.05 2.85 5.9 3.15 ;
      RECT 4.05 2.8 4.55 3.15 ;
      RECT 1.45 2.85 3.75 3.15 ;
      RECT 3.45 2.05 3.75 3.15 ;
      RECT 1.45 2.15 1.75 3.15 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 3.45 2.05 4.45 2.4 ;
      RECT 3.95 2 4.45 2.4 ;
    LAYER VIA12 ;
      RECT 5.52 2.87 5.78 3.13 ;
      RECT 4.17 2.87 4.43 3.13 ;
      RECT 4.07 2.07 4.33 2.33 ;
      RECT 2.32 3.57 2.58 3.83 ;
      RECT 1.47 2.22 1.73 2.48 ;
    LAYER MET1 ;
      RECT 4.4 3.5 4.7 5.2 ;
      RECT 2.95 3.5 5.1 3.8 ;
      RECT 4.8 1.55 5.1 3.8 ;
      RECT 2.95 2.75 3.25 3.8 ;
      RECT 2.8 2.75 3.25 3.2 ;
      RECT 4.4 1.55 5.1 1.8 ;
      RECT 4.4 0.95 4.7 1.8 ;
      RECT 2.4 3.5 2.7 5.2 ;
      RECT 2.1 1.55 2.4 3.9 ;
      RECT 2.4 0.95 2.7 1.8 ;
      RECT 1.45 0.95 1.75 5.2 ;
      RECT 1.35 2.15 1.85 2.55 ;
      RECT 5.4 2.85 5.9 3.15 ;
      RECT 4.05 2.8 4.55 3.25 ;
      RECT 3.95 2.05 4.45 2.35 ;
  END
END gf180mcu_osu_sc_gp9t3v3__lshifup

MACRO gf180mcu_osu_sc_gp9t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux2_1 0 0 ;
  SIZE 5.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.1 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.1 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 2.15 2.85 2.55 ;
        RECT 2.25 0.95 2.5 5.2 ;
      LAYER MET2 ;
        RECT 2.35 2.15 2.85 2.55 ;
      LAYER VIA12 ;
        RECT 2.47 2.22 2.73 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.25 2.15 4.75 2.55 ;
        RECT 4.25 0.95 4.5 5.2 ;
      LAYER MET2 ;
        RECT 4.25 2.15 4.75 2.55 ;
      LAYER VIA12 ;
        RECT 4.37 2.22 4.63 2.48 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 2.85 1.05 3.15 ;
      LAYER MET2 ;
        RECT 0.55 2.8 1.05 3.2 ;
      LAYER VIA12 ;
        RECT 0.67 2.87 0.93 3.13 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 4.05 3.4 4.55 ;
        RECT 3.1 0.95 3.35 5.2 ;
      LAYER MET2 ;
        RECT 3 4.1 3.5 4.5 ;
      LAYER VIA12 ;
        RECT 3.12 4.17 3.38 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 3.55 3 4.05 3.4 ;
      RECT 1.45 3 1.95 3.4 ;
      RECT 1.45 3.05 4.05 3.35 ;
    LAYER VIA12 ;
      RECT 3.67 3.07 3.93 3.33 ;
      RECT 1.57 3.07 1.83 3.33 ;
    LAYER MET1 ;
      RECT 1.4 0.95 1.65 5.2 ;
      RECT 1.4 3.05 1.95 3.35 ;
      RECT 1.4 2 2 2.3 ;
      RECT 3.65 2.9 3.95 3.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux2_1

MACRO gf180mcu_osu_sc_gp9t3v3__nand2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nand2_1 0 0 ;
  SIZE 3.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.1 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.1 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2 2.85 2.5 3.15 ;
      LAYER MET2 ;
        RECT 2 2.8 2.5 3.2 ;
      LAYER VIA12 ;
        RECT 2.12 2.87 2.38 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 1.5 1.65 5.2 ;
        RECT 0.7 1.5 1.65 1.75 ;
        RECT 0.7 0.95 0.95 1.75 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__nand2_1

MACRO gf180mcu_osu_sc_gp9t3v3__nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__nor2_1 0 0 ;
  SIZE 2.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.8 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 3.6 2.2 5.2 ;
        RECT 1.25 3.6 2.2 3.85 ;
        RECT 1.15 3.5 1.65 3.8 ;
        RECT 1.25 0.95 1.5 3.85 ;
      LAYER MET2 ;
        RECT 1.15 3.45 1.65 3.85 ;
      LAYER VIA12 ;
        RECT 1.27 3.52 1.53 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__nor2_1

MACRO gf180mcu_osu_sc_gp9t3v3__oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai21_1 0 0 ;
  SIZE 4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4 6.15 ;
        RECT 3.05 4.45 3.3 6.15 ;
        RECT 0.65 3.5 0.9 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4 0.6 ;
        RECT 1.35 0 1.6 1.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.85 2.15 3.15 ;
      LAYER MET2 ;
        RECT 1.65 2.8 2.15 3.2 ;
      LAYER VIA12 ;
        RECT 1.77 2.87 2.03 3.13 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 2.2 2.85 2.5 ;
      LAYER MET2 ;
        RECT 2.35 2.15 2.85 2.55 ;
      LAYER VIA12 ;
        RECT 2.47 2.22 2.73 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 3.5 3.5 3.8 ;
        RECT 3.1 3.45 3.45 3.8 ;
        RECT 3.15 0.95 3.4 3.8 ;
        RECT 2.1 3.5 2.45 5.2 ;
      LAYER MET2 ;
        RECT 3 3.5 3.5 3.8 ;
        RECT 3.05 3.45 3.45 3.85 ;
      LAYER VIA12 ;
        RECT 3.12 3.52 3.38 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.65 2.55 1.9 ;
      RECT 2.2 0.95 2.55 1.9 ;
      RECT 0.5 0.95 0.75 1.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai21_1

MACRO gf180mcu_osu_sc_gp9t3v3__oai22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai22_1 0 0 ;
  SIZE 5.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.5 6.15 ;
        RECT 3.6 3.5 3.85 6.15 ;
        RECT 0.65 3.5 0.9 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.5 0.6 ;
        RECT 1.35 0 1.6 1.45 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.7 2.2 1.2 2.5 ;
      LAYER MET2 ;
        RECT 0.7 2.15 1.2 2.55 ;
      LAYER VIA12 ;
        RECT 0.82 2.22 1.08 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.2 2.15 2.5 ;
      LAYER MET2 ;
        RECT 1.65 2.15 2.15 2.55 ;
      LAYER VIA12 ;
        RECT 1.77 2.22 2.03 2.48 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 2.2 3.05 2.5 ;
      LAYER MET2 ;
        RECT 2.55 2.15 3.05 2.55 ;
      LAYER VIA12 ;
        RECT 2.67 2.22 2.93 2.48 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 2.2 3.85 2.5 ;
      LAYER MET2 ;
        RECT 3.35 2.15 3.85 2.55 ;
      LAYER VIA12 ;
        RECT 3.47 2.22 3.73 2.48 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.5 0.85 5 1.15 ;
        RECT 2.1 2.75 4.9 3.05 ;
        RECT 4.6 0.85 4.9 3.05 ;
        RECT 2.1 2.75 2.45 5.2 ;
        RECT 3.05 0.85 3.55 1.2 ;
        RECT 3.15 0.85 3.4 1.45 ;
      LAYER MET2 ;
        RECT 3.05 0.85 5 1.15 ;
        RECT 4.55 0.8 4.95 1.2 ;
        RECT 3.05 0.8 3.55 1.2 ;
      LAYER VIA12 ;
        RECT 3.17 0.87 3.43 1.13 ;
        RECT 4.62 0.87 4.88 1.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.7 4.25 1.95 ;
      RECT 4 0.95 4.25 1.95 ;
      RECT 2.2 0.95 2.55 1.95 ;
      RECT 0.5 0.95 0.75 1.95 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai22_1

MACRO gf180mcu_osu_sc_gp9t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai31_1 0 0 ;
  SIZE 4.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.9 6.15 ;
        RECT 3.95 4.45 4.2 6.15 ;
        RECT 1 3.5 1.25 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.9 0.6 ;
        RECT 2.25 0 2.5 1.4 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 2.2 2.25 2.5 ;
      LAYER MET2 ;
        RECT 1.75 2.15 2.25 2.55 ;
      LAYER VIA12 ;
        RECT 1.87 2.22 2.13 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 2.85 3.05 3.15 ;
      LAYER MET2 ;
        RECT 2.55 2.8 3.05 3.2 ;
      LAYER VIA12 ;
        RECT 2.67 2.87 2.93 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 2.2 1.25 2.5 ;
      LAYER MET2 ;
        RECT 0.75 2.15 1.25 2.55 ;
      LAYER VIA12 ;
        RECT 0.87 2.22 1.13 2.48 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.25 2.2 3.75 2.5 ;
      LAYER MET2 ;
        RECT 3.25 2.15 3.75 2.55 ;
      LAYER VIA12 ;
        RECT 3.37 2.22 3.63 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 3.5 4.4 3.8 ;
        RECT 4 3.45 4.35 3.8 ;
        RECT 4.05 0.95 4.3 3.8 ;
        RECT 3 3.5 3.35 5.2 ;
      LAYER MET2 ;
        RECT 3.9 3.5 4.4 3.8 ;
        RECT 3.95 3.45 4.35 3.85 ;
      LAYER VIA12 ;
        RECT 4.02 3.52 4.28 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.65 3.45 1.9 ;
      RECT 3.1 0.95 3.45 1.9 ;
      RECT 1.4 0.95 1.65 1.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai31_1

MACRO gf180mcu_osu_sc_gp9t3v3__or2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__or2_1 0 0 ;
  SIZE 3.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.8 6.15 ;
        RECT 1.95 4.3 2.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.45 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.9 2.2 1.4 2.5 ;
      LAYER MET2 ;
        RECT 0.9 2.15 1.4 2.55 ;
      LAYER VIA12 ;
        RECT 1.02 2.22 1.28 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.85 2.15 3.15 ;
      LAYER MET2 ;
        RECT 1.65 2.8 2.15 3.2 ;
      LAYER VIA12 ;
        RECT 1.77 2.87 2.03 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 1.45 3.45 1.75 ;
        RECT 2.95 0.95 3.2 1.8 ;
        RECT 2.95 3.5 3.45 3.8 ;
        RECT 2.95 3.5 3.2 5.2 ;
      LAYER MET2 ;
        RECT 2.95 3.45 3.45 3.85 ;
        RECT 2.95 1.4 3.45 1.8 ;
        RECT 3.05 1.4 3.35 3.85 ;
      LAYER VIA12 ;
        RECT 3.07 3.52 3.33 3.78 ;
        RECT 3.07 1.47 3.33 1.73 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 2.95 0.8 5.2 ;
      RECT 0.55 3.75 2.7 4.05 ;
      RECT 2.4 2.95 2.7 4.05 ;
      RECT 2.4 2.95 2.95 3.25 ;
      RECT 0.4 1.7 0.65 3.25 ;
      RECT 0.4 1.7 1.5 1.95 ;
      RECT 1.25 0.95 1.5 1.95 ;
  END
END gf180mcu_osu_sc_gp9t3v3__or2_1

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_1 0 0 ;
  SIZE 4.15 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.15 6.15 ;
        RECT 2.35 3.9 2.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.15 0.6 ;
        RECT 2.35 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.85 2.45 3.15 ;
        RECT 2 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.2 3.5 3.7 3.8 ;
        RECT 3.4 1.5 3.65 3.8 ;
        RECT 3.3 3.4 3.55 5.2 ;
        RECT 3.3 0.95 3.55 1.8 ;
      LAYER MET2 ;
        RECT 3.2 3.45 3.7 3.85 ;
      LAYER VIA12 ;
        RECT 3.32 3.52 3.58 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.95 3.4 1.2 5.2 ;
      RECT 0.95 3.4 2.95 3.65 ;
      RECT 2.7 2.15 2.95 3.65 ;
      RECT 1.65 2.15 3.15 2.45 ;
      RECT 1.65 1.55 1.9 2.45 ;
      RECT 0.95 1.55 1.9 1.8 ;
      RECT 0.95 0.95 1.2 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_1

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_16 0 0 ;
  SIZE 16.85 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 16.85 6.15 ;
        RECT 16.05 3.5 16.3 6.15 ;
        RECT 14.35 3.5 14.6 6.15 ;
        RECT 12.65 3.5 12.9 6.15 ;
        RECT 10.95 3.5 11.2 6.15 ;
        RECT 9.25 3.5 9.5 6.15 ;
        RECT 7.55 3.5 7.8 6.15 ;
        RECT 5.85 3.5 6.1 6.15 ;
        RECT 4.15 3.5 4.4 6.15 ;
        RECT 2.35 3.9 2.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 16.85 0.6 ;
        RECT 16.05 0 16.3 1.8 ;
        RECT 14.35 0 14.6 1.8 ;
        RECT 12.65 0 12.9 1.8 ;
        RECT 10.95 0 11.2 1.8 ;
        RECT 9.25 0 9.5 1.8 ;
        RECT 7.55 0 7.8 1.8 ;
        RECT 5.85 0 6.1 1.8 ;
        RECT 4.15 0 4.4 1.8 ;
        RECT 2.35 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.85 2.45 3.15 ;
        RECT 2 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.1 3.5 15.6 3.8 ;
        RECT 15.2 0.95 15.45 5.2 ;
        RECT 3.3 2.95 15.45 3.25 ;
        RECT 3.3 2.05 15.45 2.35 ;
        RECT 13.5 0.95 13.75 5.2 ;
        RECT 11.8 0.95 12.05 5.2 ;
        RECT 10.1 0.95 10.35 5.2 ;
        RECT 8.4 0.95 8.65 5.2 ;
        RECT 6.7 0.95 6.95 5.2 ;
        RECT 5 0.95 5.25 5.2 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 15.1 3.45 15.6 3.85 ;
      LAYER VIA12 ;
        RECT 15.22 3.52 15.48 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.95 3.4 1.2 5.2 ;
      RECT 0.95 3.4 2.95 3.65 ;
      RECT 2.7 2.05 2.95 3.65 ;
      RECT 2.7 2.05 3.05 2.55 ;
      RECT 1.65 2.15 3.05 2.45 ;
      RECT 1.65 1.55 1.9 2.45 ;
      RECT 0.95 1.55 1.9 1.8 ;
      RECT 0.95 0.95 1.2 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_16

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_2 0 0 ;
  SIZE 4.95 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.95 6.15 ;
        RECT 4.15 3.5 4.4 6.15 ;
        RECT 2.35 3.9 2.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.95 0.6 ;
        RECT 4.15 0 4.4 1.8 ;
        RECT 2.35 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.85 2.45 3.15 ;
        RECT 2 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.2 3.5 3.7 3.8 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 3.2 3.45 3.7 3.85 ;
      LAYER VIA12 ;
        RECT 3.32 3.52 3.58 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.95 3.4 1.2 5.2 ;
      RECT 0.95 3.4 2.95 3.65 ;
      RECT 2.7 2.05 2.95 3.65 ;
      RECT 2.7 2.05 3.05 2.55 ;
      RECT 1.65 2.15 3.05 2.45 ;
      RECT 1.65 1.55 1.9 2.45 ;
      RECT 0.95 1.55 1.9 1.8 ;
      RECT 0.95 0.95 1.2 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_2

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_4 0 0 ;
  SIZE 6.7 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 6.7 6.15 ;
        RECT 5.85 3.5 6.1 6.15 ;
        RECT 4.15 3.5 4.4 6.15 ;
        RECT 2.35 3.9 2.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.7 0.6 ;
        RECT 5.85 0 6.1 1.8 ;
        RECT 4.15 0 4.4 1.8 ;
        RECT 2.35 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.85 2.45 3.15 ;
        RECT 2 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.9 3.5 5.4 3.8 ;
        RECT 5 0.95 5.25 5.2 ;
        RECT 3.3 2.95 5.25 3.25 ;
        RECT 3.3 2.05 5.25 2.35 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 4.9 3.45 5.4 3.85 ;
      LAYER VIA12 ;
        RECT 5.02 3.52 5.28 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.95 3.4 1.2 5.2 ;
      RECT 0.95 3.4 2.95 3.65 ;
      RECT 2.7 2.05 2.95 3.65 ;
      RECT 2.7 2.05 3.05 2.55 ;
      RECT 1.65 2.15 3.05 2.45 ;
      RECT 1.65 1.55 1.9 2.45 ;
      RECT 0.95 1.55 1.9 1.8 ;
      RECT 0.95 0.95 1.2 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_4

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_8 0 0 ;
  SIZE 10.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 10.1 6.15 ;
        RECT 9.25 3.5 9.5 6.15 ;
        RECT 7.55 3.5 7.8 6.15 ;
        RECT 5.85 3.5 6.1 6.15 ;
        RECT 4.15 3.5 4.4 6.15 ;
        RECT 2.35 3.9 2.7 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 10.1 0.6 ;
        RECT 9.25 0 9.5 1.8 ;
        RECT 7.55 0 7.8 1.8 ;
        RECT 5.85 0 6.1 1.8 ;
        RECT 4.15 0 4.4 1.8 ;
        RECT 2.35 0 2.7 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 2.85 2.45 3.15 ;
      LAYER MET2 ;
        RECT 1.95 2.85 2.45 3.15 ;
        RECT 2 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.07 2.87 2.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.3 3.5 8.8 3.8 ;
        RECT 8.4 0.95 8.65 5.2 ;
        RECT 3.3 2.95 8.65 3.25 ;
        RECT 3.3 2.05 8.65 2.35 ;
        RECT 6.7 0.95 6.95 5.2 ;
        RECT 5 0.95 5.25 5.2 ;
        RECT 3.3 0.95 3.55 5.2 ;
      LAYER MET2 ;
        RECT 8.3 3.45 8.8 3.85 ;
      LAYER VIA12 ;
        RECT 8.42 3.52 8.68 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.95 3.4 1.2 5.2 ;
      RECT 0.95 3.4 2.95 3.65 ;
      RECT 2.7 2.05 2.95 3.65 ;
      RECT 2.7 2.05 3.05 2.55 ;
      RECT 1.65 2.15 3.05 2.45 ;
      RECT 1.65 1.55 1.9 2.45 ;
      RECT 0.95 1.55 1.9 1.8 ;
      RECT 0.95 0.95 1.2 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_8

MACRO gf180mcu_osu_sc_gp9t3v3__tiehi
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tiehi 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 3.5 1.8 3.8 ;
        RECT 1.4 3.45 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.3 3.45 1.8 3.85 ;
      LAYER VIA12 ;
        RECT 1.42 3.52 1.68 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.15 2.2 1.65 2.45 ;
      RECT 1.4 0.95 1.65 2.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tiehi

MACRO gf180mcu_osu_sc_gp9t3v3__tielo
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tielo 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 1.55 1.8 1.85 ;
        RECT 1.4 0.95 1.65 1.9 ;
      LAYER MET2 ;
        RECT 1.3 1.5 1.8 1.9 ;
      LAYER VIA12 ;
        RECT 1.42 1.57 1.68 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 2.9 1.65 5.2 ;
      RECT 1.15 2.9 1.65 3.15 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tielo

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_1 0 0 ;
  SIZE 3.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.5 6.15 ;
        RECT 1.15 3.5 1.4 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.5 0.6 ;
        RECT 1.15 0 1.4 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.15 2.1 2.45 2.6 ;
      LAYER MET2 ;
        RECT 2.05 2.15 2.55 2.55 ;
      LAYER VIA12 ;
        RECT 2.17 2.22 2.43 2.48 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.5 2.2 1 2.5 ;
      LAYER MET2 ;
        RECT 0.5 2.15 1 2.55 ;
      LAYER VIA12 ;
        RECT 0.62 2.22 0.88 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.2 2.85 1.7 3.15 ;
      LAYER MET2 ;
        RECT 1.2 2.8 1.7 3.2 ;
      LAYER VIA12 ;
        RECT 1.32 2.87 1.58 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.45 3.5 2.95 3.8 ;
        RECT 2.7 1.55 2.95 3.8 ;
        RECT 2.55 3.4 2.8 5.2 ;
        RECT 2.55 0.95 2.8 1.8 ;
      LAYER MET2 ;
        RECT 2.45 3.45 2.95 3.85 ;
      LAYER VIA12 ;
        RECT 2.57 3.52 2.83 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__tinv_1

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_16 0 0 ;
  SIZE 18.3 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 18.3 6.15 ;
        RECT 17.45 3.5 17.7 6.15 ;
        RECT 15.75 3.5 16 6.15 ;
        RECT 14.05 3.5 14.3 6.15 ;
        RECT 12.35 3.5 12.6 6.15 ;
        RECT 10.65 3.5 10.9 6.15 ;
        RECT 8.95 3.5 9.2 6.15 ;
        RECT 7.25 3.5 7.5 6.15 ;
        RECT 5.55 3.5 5.8 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 1.1 3.5 1.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 18.3 0.6 ;
        RECT 17.45 0 17.7 1.8 ;
        RECT 15.75 0 16 1.8 ;
        RECT 14.05 0 14.3 1.8 ;
        RECT 12.35 0 12.6 1.8 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.95 0 9.2 1.8 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.1 0 1.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 1.45 2.25 2.9 ;
      LAYER MET2 ;
        RECT 1.85 1.5 2.35 1.9 ;
      LAYER VIA12 ;
        RECT 1.97 1.57 2.23 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.6 3.5 17.15 3.8 ;
        RECT 16.6 0.95 16.85 5.2 ;
        RECT 4.7 3 16.85 3.25 ;
        RECT 4.7 2.05 16.85 2.3 ;
        RECT 14.9 0.95 15.15 5.2 ;
        RECT 13.2 0.95 13.45 5.2 ;
        RECT 11.5 0.95 11.75 5.2 ;
        RECT 9.8 0.95 10.05 5.2 ;
        RECT 8.1 0.95 8.35 5.2 ;
        RECT 6.4 0.95 6.65 5.2 ;
        RECT 4.7 0.95 4.95 5.2 ;
      LAYER MET2 ;
        RECT 16.65 3.5 17.15 3.8 ;
        RECT 16.7 3.45 17.1 3.85 ;
      LAYER VIA12 ;
        RECT 16.77 3.52 17.03 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.4 2.8 3.95 3.2 ;
    LAYER VIA12 ;
      RECT 3.57 2.87 3.83 3.13 ;
      RECT 2.52 2.87 2.78 3.13 ;
    LAYER MET1 ;
      RECT 3 3.5 3.25 5.2 ;
      RECT 3.05 2.2 3.3 3.7 ;
      RECT 4.15 2.1 4.4 2.55 ;
      RECT 3 0.95 3.25 2.55 ;
      RECT 3 2.2 4.4 2.45 ;
      RECT 2.5 0.95 2.75 5.2 ;
      RECT 2.5 2.75 2.8 3.25 ;
      RECT 3.55 2.75 3.85 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_16

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_2
  CLASS CORE ;
  ORIGIN 3.3 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_2 -3.3 0 ;
  SIZE 6.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -3.3 5.55 3.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
        RECT -2.2 3.5 -1.95 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -3.3 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
        RECT -2.2 0 -1.95 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -1.35 1.45 -1.05 2.9 ;
      LAYER MET2 ;
        RECT -1.45 1.5 -0.95 1.9 ;
      LAYER VIA12 ;
        RECT -1.33 1.57 -1.07 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -2.85 2.2 -2.35 2.5 ;
      LAYER MET2 ;
        RECT -2.85 2.15 -2.35 2.55 ;
      LAYER VIA12 ;
        RECT -2.73 2.22 -2.47 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -2.15 2.85 -1.65 3.15 ;
      LAYER MET2 ;
        RECT -2.15 2.8 -1.65 3.2 ;
      LAYER VIA12 ;
        RECT -2.03 2.87 -1.77 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 3 2.65 3.25 ;
        RECT 2.4 2.05 2.65 3.25 ;
        RECT 1.4 2.05 2.65 2.3 ;
        RECT 1.4 3 1.95 3.9 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.55 3.5 2.05 3.8 ;
        RECT 1.6 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.67 3.52 1.93 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT -0.9 2.8 0.65 3.2 ;
    LAYER VIA12 ;
      RECT 0.27 2.87 0.53 3.13 ;
      RECT -0.78 2.87 -0.52 3.13 ;
    LAYER MET1 ;
      RECT -0.3 3.5 -0.05 5.2 ;
      RECT -0.25 2.2 0 3.7 ;
      RECT 0.85 2.1 1.1 2.55 ;
      RECT -0.3 0.95 -0.05 2.55 ;
      RECT -0.3 2.2 1.1 2.45 ;
      RECT -0.8 0.95 -0.55 5.2 ;
      RECT -0.8 2.75 -0.5 3.25 ;
      RECT 0.25 2.75 0.55 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_2

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_4 0 0 ;
  SIZE 8.1 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.1 6.15 ;
        RECT 7.3 3.5 7.55 6.15 ;
        RECT 5.55 3.5 5.8 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 1.1 3.5 1.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.1 0.6 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.1 0 1.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 1.45 2.25 2.9 ;
      LAYER MET2 ;
        RECT 1.85 1.5 2.35 1.9 ;
      LAYER VIA12 ;
        RECT 1.97 1.57 2.23 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.4 3.5 7.05 3.8 ;
        RECT 6.4 0.95 6.65 5.2 ;
        RECT 4.7 3 6.65 3.25 ;
        RECT 4.7 2.05 6.65 2.3 ;
        RECT 4.7 0.95 4.95 5.2 ;
      LAYER MET2 ;
        RECT 6.55 3.5 7.05 3.8 ;
        RECT 6.6 3.45 7 3.85 ;
      LAYER VIA12 ;
        RECT 6.67 3.52 6.93 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.4 2.8 3.95 3.2 ;
    LAYER VIA12 ;
      RECT 3.57 2.87 3.83 3.13 ;
      RECT 2.52 2.87 2.78 3.13 ;
    LAYER MET1 ;
      RECT 3 3.5 3.25 5.2 ;
      RECT 3.05 2.2 3.3 3.7 ;
      RECT 4.15 2.1 4.4 2.55 ;
      RECT 3 0.95 3.25 2.55 ;
      RECT 3 2.2 4.4 2.45 ;
      RECT 2.5 0.95 2.75 5.2 ;
      RECT 2.5 2.75 2.8 3.25 ;
      RECT 3.55 2.75 3.85 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_4

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_8 0 0 ;
  SIZE 11.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 11.5 6.15 ;
        RECT 10.7 3.5 10.95 6.15 ;
        RECT 8.95 3.5 9.2 6.15 ;
        RECT 7.25 3.5 7.5 6.15 ;
        RECT 5.55 3.5 5.8 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 1.1 3.5 1.35 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 11.5 0.6 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.95 0 9.2 1.8 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 5.55 0 5.8 1.8 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.1 0 1.35 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 1.45 2.25 2.9 ;
      LAYER MET2 ;
        RECT 1.85 1.5 2.35 1.9 ;
      LAYER VIA12 ;
        RECT 1.97 1.57 2.23 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 2.2 0.95 2.5 ;
      LAYER MET2 ;
        RECT 0.45 2.15 0.95 2.55 ;
      LAYER VIA12 ;
        RECT 0.57 2.22 0.83 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.15 2.85 1.65 3.15 ;
      LAYER MET2 ;
        RECT 1.15 2.8 1.65 3.2 ;
      LAYER VIA12 ;
        RECT 1.27 2.87 1.53 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.8 3.5 10.45 3.8 ;
        RECT 9.8 0.95 10.05 5.2 ;
        RECT 4.7 3 10.05 3.25 ;
        RECT 4.7 2.05 10.05 2.3 ;
        RECT 8.1 0.95 8.35 5.2 ;
        RECT 6.4 0.95 6.65 5.2 ;
        RECT 4.7 0.95 4.95 5.2 ;
      LAYER MET2 ;
        RECT 9.95 3.5 10.45 3.8 ;
        RECT 10 3.45 10.4 3.85 ;
      LAYER VIA12 ;
        RECT 10.07 3.52 10.33 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.4 2.8 3.95 3.2 ;
    LAYER VIA12 ;
      RECT 3.57 2.87 3.83 3.13 ;
      RECT 2.52 2.87 2.78 3.13 ;
    LAYER MET1 ;
      RECT 3 3.5 3.25 5.2 ;
      RECT 3.05 2.2 3.3 3.7 ;
      RECT 4.15 2.1 4.4 2.55 ;
      RECT 3 0.95 3.25 2.55 ;
      RECT 3 2.2 4.4 2.45 ;
      RECT 2.5 0.95 2.75 5.2 ;
      RECT 2.5 2.75 2.8 3.25 ;
      RECT 3.55 2.75 3.85 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_8

MACRO gf180mcu_osu_sc_gp9t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xnor2_1 0 0 ;
  SIZE 6.4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 6.4 6.15 ;
        RECT 4.7 4.6 4.95 6.15 ;
        RECT 1.4 4.6 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.4 0.6 ;
        RECT 4.7 0 4.95 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.5 3 4 3.3 ;
        RECT 1.25 2.2 1.75 2.5 ;
      LAYER MET2 ;
        RECT 3.55 2.95 4 3.35 ;
        RECT 3.7 0.9 4 3.35 ;
        RECT 3.6 2.9 3.95 3.4 ;
        RECT 1.35 0.9 4 1.2 ;
        RECT 1.3 2.15 1.7 2.55 ;
        RECT 1.35 0.9 1.65 2.6 ;
      LAYER VIA12 ;
        RECT 1.37 2.22 1.63 2.48 ;
        RECT 3.62 3.02 3.88 3.28 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.55 2.2 5.05 2.5 ;
      LAYER MET2 ;
        RECT 4.55 2.2 5.05 2.5 ;
        RECT 4.6 2.15 5 2.55 ;
        RECT 4.65 2.1 4.95 2.6 ;
      LAYER VIA12 ;
        RECT 4.67 2.22 4.93 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 1.4 3.3 1.95 ;
        RECT 3.05 0.95 3.3 1.95 ;
        RECT 3.05 4.05 3.3 5.2 ;
        RECT 3 4.05 3.3 4.75 ;
      LAYER MET2 ;
        RECT 2.9 1.5 3.4 1.9 ;
        RECT 2.95 4.1 3.35 4.5 ;
        RECT 3 4.05 3.3 4.75 ;
        RECT 2.95 1.5 3.25 4.5 ;
      LAYER VIA12 ;
        RECT 3.02 4.17 3.28 4.43 ;
        RECT 3.02 1.57 3.28 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.55 0.95 5.8 5.2 ;
      RECT 2.75 3.55 5.8 3.8 ;
      RECT 2.75 2.9 3.05 3.8 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 3 2.4 3.3 ;
      RECT 2.1 2.2 2.4 3.3 ;
      RECT 2.1 2.2 3.5 2.5 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xnor2_1

MACRO gf180mcu_osu_sc_gp9t3v3__xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xor2_1 0 0 ;
  SIZE 6.7 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 6.7 6.15 ;
        RECT 5 3.8 5.25 6.15 ;
        RECT 1.4 3.8 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.7 0.6 ;
        RECT 5 0 5.25 1.75 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.1 2.2 1.6 2.5 ;
      LAYER MET2 ;
        RECT 1.1 2.2 1.6 2.5 ;
        RECT 1.15 2.15 1.55 2.55 ;
      LAYER VIA12 ;
        RECT 1.22 2.22 1.48 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.1 2.2 5.6 2.5 ;
        RECT 2.35 2 5.45 2.3 ;
      LAYER MET2 ;
        RECT 5.1 2.2 5.6 2.5 ;
        RECT 5.15 2.15 5.55 2.55 ;
      LAYER VIA12 ;
        RECT 5.22 2.22 5.48 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.05 1.4 3.55 1.7 ;
        RECT 3.15 1.3 3.45 1.75 ;
        RECT 3.2 0.95 3.45 1.75 ;
        RECT 3.05 4.15 3.55 4.45 ;
        RECT 3.2 4.15 3.45 5.2 ;
        RECT 3.15 4.15 3.45 4.55 ;
      LAYER MET2 ;
        RECT 3.05 1.35 3.55 1.75 ;
        RECT 3.1 4.1 3.5 4.5 ;
        RECT 3.15 1.35 3.45 4.55 ;
      LAYER VIA12 ;
        RECT 3.17 4.17 3.43 4.43 ;
        RECT 3.17 1.42 3.43 1.68 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.85 0.95 6.1 5.2 ;
      RECT 2.7 3.65 4.7 3.9 ;
      RECT 4.45 2.55 4.7 3.9 ;
      RECT 2.7 3.05 3 3.9 ;
      RECT 4.45 3.1 6.1 3.4 ;
      RECT 2.6 3.05 3.1 3.3 ;
      RECT 4.45 2.55 4.75 3.4 ;
      RECT 4.35 2.55 4.85 2.85 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 3.65 2.55 3.95 3.4 ;
      RECT 0.55 3 2.35 3.25 ;
      RECT 2.05 2.55 2.35 3.25 ;
      RECT 2.05 2.55 3.95 2.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xor2_1

END LIBRARY
