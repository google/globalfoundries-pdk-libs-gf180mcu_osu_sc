magic
tech gf180mcuC
timestamp 1660080223
<< nwell >>
rect 0 97 76 159
<< nmos >>
rect 16 16 22 33
rect 33 16 39 33
rect 50 16 56 33
<< pmos >>
rect 19 106 25 140
rect 30 106 36 140
rect 50 106 56 140
<< ndiff >>
rect 6 31 16 33
rect 6 18 8 31
rect 13 18 16 31
rect 6 16 16 18
rect 22 31 33 33
rect 22 18 25 31
rect 30 18 33 31
rect 22 16 33 18
rect 39 31 50 33
rect 39 18 42 31
rect 47 18 50 31
rect 39 16 50 18
rect 56 31 66 33
rect 56 18 59 31
rect 64 18 66 31
rect 56 16 66 18
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 106 30 140
rect 36 138 50 140
rect 36 108 39 138
rect 47 108 50 138
rect 36 106 50 108
rect 56 138 66 140
rect 56 108 59 138
rect 64 108 66 138
rect 56 106 66 108
<< ndiffc >>
rect 8 18 13 31
rect 25 18 30 31
rect 42 18 47 31
rect 59 18 64 31
<< pdiffc >>
rect 11 108 16 138
rect 39 108 47 138
rect 59 108 64 138
<< psubdiff >>
rect 9 7 18 9
rect 9 2 11 7
rect 16 2 18 7
rect 9 0 18 2
rect 33 7 42 9
rect 33 2 35 7
rect 40 2 42 7
rect 33 0 42 2
rect 57 7 66 9
rect 57 2 59 7
rect 64 2 66 7
rect 57 0 66 2
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
<< psubdiffcont >>
rect 11 2 16 7
rect 35 2 40 7
rect 59 2 64 7
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
<< polysilicon >>
rect 19 140 25 145
rect 30 140 36 145
rect 50 140 56 145
rect 19 102 25 106
rect 16 97 25 102
rect 30 103 36 106
rect 30 97 39 103
rect 16 75 22 97
rect 16 73 28 75
rect 16 67 20 73
rect 26 67 28 73
rect 16 65 28 67
rect 16 33 22 65
rect 33 62 39 97
rect 50 88 56 106
rect 44 86 56 88
rect 44 80 46 86
rect 52 80 56 86
rect 44 78 56 80
rect 33 60 43 62
rect 33 54 35 60
rect 41 54 43 60
rect 33 52 43 54
rect 33 33 39 52
rect 50 33 56 78
rect 16 11 22 16
rect 33 11 39 16
rect 50 11 56 16
<< polycontact >>
rect 20 67 26 73
rect 46 80 52 86
rect 35 54 41 60
<< metal1 >>
rect 0 154 76 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 76 154
rect 0 147 76 148
rect 11 138 16 140
rect 11 107 16 108
rect 8 102 16 107
rect 39 138 47 147
rect 39 106 47 108
rect 59 138 64 140
rect 8 86 13 102
rect 59 99 64 108
rect 59 93 61 99
rect 67 93 69 99
rect 8 80 46 86
rect 52 80 54 86
rect 8 46 13 80
rect 18 67 20 73
rect 26 67 28 73
rect 33 54 35 60
rect 41 54 43 60
rect 8 41 30 46
rect 8 31 13 33
rect 8 9 13 18
rect 25 31 30 41
rect 25 16 30 18
rect 42 31 47 33
rect 42 9 47 18
rect 59 31 64 93
rect 59 16 64 18
rect 0 8 76 9
rect 0 2 11 8
rect 17 2 35 8
rect 41 2 59 8
rect 65 2 76 8
rect 0 -3 76 2
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 61 93 67 99
rect 46 80 52 86
rect 20 67 26 73
rect 35 54 41 60
rect 11 7 17 8
rect 11 2 16 7
rect 16 2 17 7
rect 35 7 41 8
rect 35 2 40 7
rect 40 2 41 7
rect 59 7 65 8
rect 59 2 64 7
rect 64 2 65 7
<< metal2 >>
rect 9 154 19 155
rect 9 148 11 154
rect 17 148 19 154
rect 9 147 19 148
rect 33 154 43 155
rect 33 148 35 154
rect 41 148 43 154
rect 33 147 43 148
rect 57 154 67 155
rect 57 148 59 154
rect 65 148 67 154
rect 57 147 67 148
rect 59 99 69 100
rect 59 93 61 99
rect 67 93 69 99
rect 59 92 69 93
rect 44 86 54 87
rect 44 80 46 86
rect 52 80 54 86
rect 44 79 54 80
rect 18 73 28 74
rect 18 67 20 73
rect 26 67 28 73
rect 18 66 28 67
rect 33 60 43 61
rect 33 54 35 60
rect 41 54 43 60
rect 33 53 43 54
rect 9 8 19 9
rect 9 2 11 8
rect 17 2 19 8
rect 9 1 19 2
rect 33 8 43 9
rect 33 2 35 8
rect 41 2 43 8
rect 33 1 43 2
rect 57 8 67 9
rect 57 2 59 8
rect 65 2 67 8
rect 57 1 67 2
<< labels >>
rlabel metal2 23 70 23 70 1 A
port 2 n
rlabel metal2 64 96 64 96 1 Y
port 3 n
rlabel metal2 14 5 14 5 1 GND
rlabel metal2 14 152 14 152 1 VDD
rlabel metal2 38 57 38 57 1 B
port 1 n
<< end >>
