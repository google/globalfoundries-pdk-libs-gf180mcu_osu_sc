# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_16 0 0 ;
  SIZE 15 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 15 6.15 ;
        RECT 14.15 3.5 14.4 6.15 ;
        RECT 12.45 3.5 12.7 6.15 ;
        RECT 10.75 3.5 11 6.15 ;
        RECT 9.05 3.5 9.3 6.15 ;
        RECT 7.35 3.5 7.6 6.15 ;
        RECT 5.65 3.5 5.9 6.15 ;
        RECT 3.95 3.5 4.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15 0.6 ;
        RECT 14.15 0 14.4 1.8 ;
        RECT 12.45 0 12.7 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 9.05 0 9.3 1.8 ;
        RECT 7.35 0 7.6 1.8 ;
        RECT 5.65 0 5.9 1.8 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.3 3.5 13.85 3.8 ;
        RECT 13.3 0.95 13.55 5.2 ;
        RECT 1.4 3 13.55 3.25 ;
        RECT 1.4 2.05 13.55 2.3 ;
        RECT 11.6 0.95 11.85 5.2 ;
        RECT 9.9 0.95 10.15 5.2 ;
        RECT 8.2 0.95 8.45 5.2 ;
        RECT 6.5 0.95 6.75 5.2 ;
        RECT 4.8 0.95 5.05 5.2 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 13.35 3.5 13.85 3.8 ;
        RECT 13.4 3.45 13.8 3.85 ;
      LAYER VIA12 ;
        RECT 13.47 3.52 13.73 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_16
