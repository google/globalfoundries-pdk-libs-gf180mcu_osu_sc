# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__clkinv_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkinv_16 0 0 ;
  SIZE 15 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 15 6.35 ;
        RECT 14.15 3.6 14.4 6.35 ;
        RECT 12.45 3.6 12.7 6.35 ;
        RECT 10.75 3.6 11 6.35 ;
        RECT 9.05 3.6 9.3 6.35 ;
        RECT 7.35 3.6 7.6 6.35 ;
        RECT 5.65 3.6 5.9 6.35 ;
        RECT 3.95 3.6 4.2 6.35 ;
        RECT 2.25 3.6 2.5 6.35 ;
        RECT 0.55 3.6 0.8 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15 0.7 ;
        RECT 14.15 0 14.4 1.9 ;
        RECT 12.45 0 12.7 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 9.05 0 9.3 1.9 ;
        RECT 7.35 0 7.6 1.9 ;
        RECT 5.65 0 5.9 1.9 ;
        RECT 3.95 0 4.2 1.9 ;
        RECT 2.25 0 2.5 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.4 2.3 0.9 2.6 ;
      LAYER Metal2 ;
        RECT 0.4 2.25 0.9 2.65 ;
      LAYER Via1 ;
        RECT 0.52 2.32 0.78 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.3 3.6 13.85 3.9 ;
        RECT 13.3 1.05 13.55 5.3 ;
        RECT 1.4 3.1 13.55 3.35 ;
        RECT 1.4 2.15 13.55 2.4 ;
        RECT 11.6 1.05 11.85 5.3 ;
        RECT 9.9 1.05 10.15 5.3 ;
        RECT 8.2 1.05 8.45 5.3 ;
        RECT 6.5 1.05 6.75 5.3 ;
        RECT 4.8 1.05 5.05 5.3 ;
        RECT 3.1 1.05 3.35 5.3 ;
        RECT 1.4 1.05 1.65 5.3 ;
      LAYER Metal2 ;
        RECT 13.35 3.6 13.85 3.9 ;
        RECT 13.4 3.55 13.8 3.95 ;
      LAYER Via1 ;
        RECT 13.47 3.62 13.73 3.88 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__clkinv_16
