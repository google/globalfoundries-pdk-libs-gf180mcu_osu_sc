* NGSPICE file created from gf180mcu_osu_sc_12T_and2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y a_12_16# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 VDD B a_12_16# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_12_16# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Y a_12_16# GND GND nmos_3p3 w=0.85u l=0.3u
X4 a_28_16# A a_12_16# GND nmos_3p3 w=0.85u l=0.3u
X5 GND B a_28_16# GND nmos_3p3 w=0.85u l=0.3u
