* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addf_1 A B CI S CO VDD VSS
X0 S a_161_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD CI a_195_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_195_21# B a_178_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_76_111# B a_59_21# VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD A a_76_111# VDD pfet_03p3 w=1.7u l=0.3u
X5 a_178_21# A a_161_21# VSS nfet_03p3 w=0.85u l=0.3u
X6 a_59_21# CI a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X7 a_9_111# B VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 a_110_21# CI VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 VDD A a_9_111# VDD pfet_03p3 w=1.7u l=0.3u
X10 a_59_21# CI a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS B a_110_21# VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS A a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X13 CO a_59_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS CI a_195_21# VSS nfet_03p3 w=0.85u l=0.3u
X15 CO a_59_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X16 VSS A a_76_21# VSS nfet_03p3 w=0.85u l=0.3u
X17 a_161_21# a_59_21# a_110_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 a_76_21# B a_59_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 a_178_111# A a_161_21# VDD pfet_03p3 w=1.7u l=0.3u
X20 a_195_111# B a_178_111# VDD pfet_03p3 w=1.7u l=0.3u
X21 a_9_21# B VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 a_110_21# A VSS VSS nfet_03p3 w=0.85u l=0.3u
X23 a_161_21# a_59_21# a_110_111# VDD pfet_03p3 w=1.7u l=0.3u
X24 a_110_111# CI VDD VDD pfet_03p3 w=1.7u l=0.3u
X25 VDD B a_110_111# VDD pfet_03p3 w=1.7u l=0.3u
X26 a_110_111# A VDD VDD pfet_03p3 w=1.7u l=0.3u
X27 S a_161_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends
