magic
tech gf180mcuC
timestamp 1659394601
<< nwell >>
rect 0 97 704 159
<< metal1 >>
rect 0 147 704 159
rect 0 -3 704 9
<< end >>
