# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_dffsr_1
  CLASS CORE ;
  ORIGIN 4.05 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_dffsr_1 -4.05 -0.15 ;
  SIZE 18.7 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.65 4 8.15 4.3 ;
        RECT 5.5 4 6.55 4.3 ;
        RECT 5.4 2 5.9 2.3 ;
        RECT 5.5 2 5.8 4.3 ;
        RECT 2.6 4 3.75 4.3 ;
        RECT 3.25 2.05 3.75 2.35 ;
        RECT 3.35 2.05 3.65 4.3 ;
      LAYER MET2 ;
        RECT 3.25 4 8.15 4.3 ;
        RECT 7.7 3.95 8.1 4.35 ;
        RECT 6.05 3.95 6.55 4.35 ;
        RECT 3.25 3.95 3.7 4.35 ;
      LAYER VIA12 ;
        RECT 3.37 4.02 3.63 4.28 ;
        RECT 6.17 4.02 6.43 4.28 ;
        RECT 7.77 4.02 8.03 4.28 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.35 2.4 3.65 ;
      LAYER MET2 ;
        RECT 1.9 3.3 2.4 3.7 ;
      LAYER VIA12 ;
        RECT 2.02 3.37 2.28 3.63 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.85 4.65 14.35 5 ;
        RECT 13.85 4.6 14.3 5 ;
        RECT 13.85 0.8 14.1 7 ;
      LAYER MET2 ;
        RECT 13.85 4.65 14.35 4.95 ;
        RECT 13.9 4.6 14.3 5 ;
      LAYER VIA12 ;
        RECT 13.97 4.67 14.23 4.93 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.15 4 13.6 4.3 ;
        RECT 13.25 1.9 13.5 4.3 ;
        RECT 12.15 1.9 13.5 2.15 ;
        RECT 12.15 4 12.4 7 ;
        RECT 12.15 0.8 12.4 2.15 ;
      LAYER MET2 ;
        RECT 13.1 4 13.6 4.3 ;
        RECT 13.15 3.95 13.55 4.35 ;
      LAYER VIA12 ;
        RECT 13.22 4.02 13.48 4.28 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -3.5 4.65 -3 4.95 ;
      LAYER MET2 ;
        RECT -3.5 4.6 -3 5 ;
      LAYER VIA12 ;
        RECT -3.38 4.67 -3.12 4.93 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.9 4 10.4 4.3 ;
        RECT -0.65 4 -0.15 4.3 ;
      LAYER MET2 ;
        RECT 9.9 3.95 10.4 4.35 ;
        RECT -0.55 5.3 10.3 5.6 ;
        RECT 10 3.95 10.3 5.6 ;
        RECT -0.65 3.95 -0.15 4.35 ;
        RECT -0.55 3.95 -0.25 5.6 ;
      LAYER VIA12 ;
        RECT -0.53 4.02 -0.27 4.28 ;
        RECT 10.02 4.02 10.28 4.28 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -4.05 7.35 14.65 7.95 ;
        RECT 13 5.3 13.25 7.95 ;
        RECT 9.7 6.55 9.95 7.95 ;
        RECT 7.25 6.05 7.5 7.95 ;
        RECT 4.45 5.3 4.7 7.95 ;
        RECT 1.4 5.3 1.65 7.95 ;
        RECT -0.2 6.05 0.05 7.95 ;
        RECT -3.5 5.3 -3.25 7.95 ;
      LAYER MET2 ;
        RECT 13.2 7.4 13.7 7.7 ;
        RECT 13.25 7.35 13.65 7.75 ;
        RECT 12 7.4 12.5 7.7 ;
        RECT 12.05 7.35 12.45 7.75 ;
        RECT 10.8 7.4 11.3 7.7 ;
        RECT 10.85 7.35 11.25 7.75 ;
        RECT 9.6 7.4 10.1 7.7 ;
        RECT 9.65 7.35 10.05 7.75 ;
        RECT 8.4 7.4 8.9 7.7 ;
        RECT 8.45 7.35 8.85 7.75 ;
        RECT 7.2 7.4 7.7 7.7 ;
        RECT 7.25 7.35 7.65 7.75 ;
        RECT 6 7.4 6.5 7.7 ;
        RECT 6.05 7.35 6.45 7.75 ;
        RECT 4.8 7.4 5.3 7.7 ;
        RECT 4.85 7.35 5.25 7.75 ;
        RECT 3.6 7.4 4.1 7.7 ;
        RECT 3.65 7.35 4.05 7.75 ;
        RECT 2.4 7.4 2.9 7.7 ;
        RECT 2.45 7.35 2.85 7.75 ;
        RECT 1.2 7.4 1.7 7.7 ;
        RECT 1.25 7.35 1.65 7.75 ;
        RECT 0 7.4 0.5 7.7 ;
        RECT 0.05 7.35 0.45 7.75 ;
        RECT -1.2 7.4 -0.7 7.7 ;
        RECT -1.15 7.35 -0.75 7.75 ;
        RECT -2.4 7.4 -1.9 7.7 ;
        RECT -2.35 7.35 -1.95 7.75 ;
        RECT -3.6 7.4 -3.1 7.7 ;
        RECT -3.55 7.35 -3.15 7.75 ;
      LAYER VIA12 ;
        RECT -3.48 7.42 -3.22 7.68 ;
        RECT -2.28 7.42 -2.02 7.68 ;
        RECT -1.08 7.42 -0.82 7.68 ;
        RECT 0.12 7.42 0.38 7.68 ;
        RECT 1.32 7.42 1.58 7.68 ;
        RECT 2.52 7.42 2.78 7.68 ;
        RECT 3.72 7.42 3.98 7.68 ;
        RECT 4.92 7.42 5.18 7.68 ;
        RECT 6.12 7.42 6.38 7.68 ;
        RECT 7.32 7.42 7.58 7.68 ;
        RECT 8.52 7.42 8.78 7.68 ;
        RECT 9.72 7.42 9.98 7.68 ;
        RECT 10.92 7.42 11.18 7.68 ;
        RECT 12.12 7.42 12.38 7.68 ;
        RECT 13.32 7.42 13.58 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -4.05 -0.15 14.65 0.45 ;
        RECT 13 -0.15 13.25 1.65 ;
        RECT 11.25 -0.15 11.5 1.65 ;
        RECT 9 -0.15 9.25 1.65 ;
        RECT 7.25 -0.15 7.5 1.65 ;
        RECT 4.45 -0.15 4.7 1.25 ;
        RECT 1.4 -0.15 1.65 1.65 ;
        RECT 0.5 -0.15 0.75 1.65 ;
        RECT -1.75 -0.15 -1.5 1.65 ;
        RECT -3.5 -0.15 -3.25 1.65 ;
      LAYER MET2 ;
        RECT 13.2 0.1 13.7 0.4 ;
        RECT 13.25 0.05 13.65 0.45 ;
        RECT 12 0.1 12.5 0.4 ;
        RECT 12.05 0.05 12.45 0.45 ;
        RECT 10.8 0.1 11.3 0.4 ;
        RECT 10.85 0.05 11.25 0.45 ;
        RECT 9.6 0.1 10.1 0.4 ;
        RECT 9.65 0.05 10.05 0.45 ;
        RECT 8.4 0.1 8.9 0.4 ;
        RECT 8.45 0.05 8.85 0.45 ;
        RECT 7.2 0.1 7.7 0.4 ;
        RECT 7.25 0.05 7.65 0.45 ;
        RECT 6 0.1 6.5 0.4 ;
        RECT 6.05 0.05 6.45 0.45 ;
        RECT 4.8 0.1 5.3 0.4 ;
        RECT 4.85 0.05 5.25 0.45 ;
        RECT 3.6 0.1 4.1 0.4 ;
        RECT 3.65 0.05 4.05 0.45 ;
        RECT 2.4 0.1 2.9 0.4 ;
        RECT 2.45 0.05 2.85 0.45 ;
        RECT 1.2 0.1 1.7 0.4 ;
        RECT 1.25 0.05 1.65 0.45 ;
        RECT 0 0.1 0.5 0.4 ;
        RECT 0.05 0.05 0.45 0.45 ;
        RECT -1.2 0.1 -0.7 0.4 ;
        RECT -1.15 0.05 -0.75 0.45 ;
        RECT -2.4 0.1 -1.9 0.4 ;
        RECT -2.35 0.05 -1.95 0.45 ;
        RECT -3.6 0.1 -3.1 0.4 ;
        RECT -3.55 0.05 -3.15 0.45 ;
      LAYER VIA12 ;
        RECT -3.48 0.12 -3.22 0.38 ;
        RECT -2.28 0.12 -2.02 0.38 ;
        RECT -1.08 0.12 -0.82 0.38 ;
        RECT 0.12 0.12 0.38 0.38 ;
        RECT 1.32 0.12 1.58 0.38 ;
        RECT 2.52 0.12 2.78 0.38 ;
        RECT 3.72 0.12 3.98 0.38 ;
        RECT 4.92 0.12 5.18 0.38 ;
        RECT 6.12 0.12 6.38 0.38 ;
        RECT 7.32 0.12 7.58 0.38 ;
        RECT 8.52 0.12 8.78 0.38 ;
        RECT 9.72 0.12 9.98 0.38 ;
        RECT 10.92 0.12 11.18 0.38 ;
        RECT 12.12 0.12 12.38 0.38 ;
        RECT 13.32 0.12 13.58 0.38 ;
    END
  END VSS
  OBS
    LAYER MET2 ;
      RECT 12.4 2.65 12.8 3.05 ;
      RECT 12.05 2.7 12.85 3 ;
      RECT -1.4 3.3 -0.9 3.7 ;
      RECT -1.3 0.75 -1 3.7 ;
      RECT -2.75 2 -2.25 2.4 ;
      RECT 10.8 1.95 11.4 2.35 ;
      RECT -2.75 2.05 -1 2.35 ;
      RECT 10.8 0.75 11.1 2.35 ;
      RECT -1.3 0.75 11.1 1.05 ;
      RECT 8.9 1.95 9.4 2.35 ;
      RECT 8.9 1.4 9.3 2.35 ;
      RECT 5.8 1.35 6.2 1.75 ;
      RECT 5.75 1.4 9.3 1.7 ;
      RECT 8.95 4.6 9.35 5 ;
      RECT 6.75 4.6 7.15 5 ;
      RECT 6.7 4.65 9.4 4.95 ;
      RECT 8.05 2.65 8.45 3.05 ;
      RECT 6.1 2.65 6.5 3.05 ;
      RECT 6.05 2.7 8.55 3 ;
      RECT 6.8 3.3 7.2 3.7 ;
      RECT 6.75 3.35 7.25 3.65 ;
      RECT 4.1 2 4.5 2.4 ;
      RECT 0.35 2 0.85 2.4 ;
      RECT 0.35 2.05 4.55 2.35 ;
      RECT 11.3 4.6 11.8 5 ;
      RECT 0.35 3.3 0.85 3.7 ;
    LAYER VIA12 ;
      RECT 12.47 2.72 12.73 2.98 ;
      RECT 11.42 4.67 11.68 4.93 ;
      RECT 11.02 2.02 11.28 2.28 ;
      RECT 9.02 2.02 9.28 2.28 ;
      RECT 9.02 4.67 9.28 4.93 ;
      RECT 8.12 2.72 8.38 2.98 ;
      RECT 6.87 3.37 7.13 3.63 ;
      RECT 6.82 4.67 7.08 4.93 ;
      RECT 6.17 2.72 6.43 2.98 ;
      RECT 5.87 1.42 6.13 1.68 ;
      RECT 4.17 2.07 4.43 2.33 ;
      RECT 0.47 2.07 0.73 2.33 ;
      RECT 0.47 3.37 0.73 3.63 ;
      RECT -1.28 3.37 -1.02 3.63 ;
      RECT -2.63 2.07 -2.37 2.33 ;
    LAYER MET1 ;
      RECT 11.4 2.7 11.65 7 ;
      RECT 9 4.55 9.3 5.05 ;
      RECT 9 4.65 11.8 4.95 ;
      RECT 10.4 2.7 12.85 3 ;
      RECT 10.4 0.8 10.65 3 ;
      RECT 10.55 6.05 10.8 7 ;
      RECT 8.85 6.05 9.1 7 ;
      RECT 8.85 6.05 10.8 6.3 ;
      RECT 8.1 4.6 8.35 7 ;
      RECT 8.1 4.6 8.65 4.85 ;
      RECT 8.4 3.4 8.65 4.85 ;
      RECT 8.1 2.6 8.4 3.65 ;
      RECT 8.1 0.8 8.35 3.65 ;
      RECT 6.7 4.65 7.2 4.95 ;
      RECT 6.8 3.35 7.1 4.95 ;
      RECT 6.75 3.35 7.25 3.65 ;
      RECT 5.85 5.8 6.1 7 ;
      RECT 4.95 5.8 6.1 6.05 ;
      RECT 4.95 3.3 5.2 6.05 ;
      RECT 4.9 1.45 5.15 3.55 ;
      RECT 4.9 1.45 6.25 1.7 ;
      RECT 5.85 1.4 6.25 1.7 ;
      RECT 5.85 0.8 6.1 1.7 ;
      RECT 4.05 4.65 4.55 4.95 ;
      RECT 4.15 2.05 4.45 4.95 ;
      RECT 4.05 2.05 4.55 2.35 ;
      RECT 3.05 4.8 3.3 7 ;
      RECT 1.4 4.8 3.3 5.05 ;
      RECT 1.4 2.1 1.65 5.05 ;
      RECT 0.35 3.35 1.65 3.65 ;
      RECT 1.4 2.1 2.4 2.35 ;
      RECT 2 1.4 2.4 2.35 ;
      RECT 2 1.4 3.3 1.65 ;
      RECT 3.05 0.8 3.3 1.65 ;
      RECT 0.65 5.55 0.9 7 ;
      RECT -1.05 5.55 -0.8 7 ;
      RECT -1.05 5.55 0.9 5.8 ;
      RECT -1.9 2.35 -1.65 7 ;
      RECT -1.9 2.35 -0.65 2.6 ;
      RECT -0.9 0.8 -0.65 2.6 ;
      RECT 0.45 2 0.7 2.4 ;
      RECT -0.9 2.05 0.85 2.35 ;
      RECT -2.65 0.8 -2.4 7 ;
      RECT -2.75 2.05 -2.25 2.35 ;
      RECT -2.65 2 -2.35 2.35 ;
      RECT 10.9 2 11.4 2.3 ;
      RECT 8.9 2 9.4 2.3 ;
      RECT 6.05 2.7 6.55 3 ;
      RECT -1.4 3.35 -0.9 3.65 ;
  END
END gf180mcu_osu_sc_12T_dffsr_1
