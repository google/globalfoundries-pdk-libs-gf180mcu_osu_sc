

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_dffsr_1 D Q QN CLK RN SN
X0 a_172_70 a_139_41 a_82_14 VDD pmos_3p3 w=34 l=6
X1 a_247_47 a_25_19 a_291_70 VDD pmos_3p3 w=34 l=6
X2 GND a_41_70 a_172_19 GND nmos_3p3 w=17 l=6
X3 VDD a_41_70 a_172_70 VDD pmos_3p3 w=34 l=6
X4 GND a_247_47 a_234_19 GND nmos_3p3 w=17 l=6
X5 VDD a_247_47 a_234_70 VDD pmos_3p3 w=34 l=6
X6 a_41_70 a_25_19 GND GND nmos_3p3 w=17 l=6
X7 a_128_19 D GND GND nmos_3p3 w=17 l=6
X8 GND a_247_47 QN GND nmos_3p3 w=17 l=6
X9 a_310_19 a_211_19 GND GND nmos_3p3 w=17 l=6
X10 a_25_19 RN GND GND nmos_3p3 w=17 l=6
X11 a_128_70 D VDD VDD pmos_3p3 w=34 l=6
X12 VDD a_247_47 QN VDD pmos_3p3 w=34 l=6
X13 VDD SN a_57_70 VDD pmos_3p3 w=34 l=6
X14 a_200_19 a_41_70 GND GND nmos_3p3 w=17 l=6
X15 a_247_47 SN a_310_19 GND nmos_3p3 w=17 l=6
X16 a_25_19 RN VDD VDD pmos_3p3 w=34 l=6
X17 a_57_70 a_25_19 a_41_70 VDD pmos_3p3 w=34 l=6
X18 a_291_70 SN VDD VDD pmos_3p3 w=34 l=6
X19 a_211_19 CLK a_200_19 GND nmos_3p3 w=17 l=6
X20 a_200_70 a_41_70 VDD VDD pmos_3p3 w=34 l=6
X21 VDD a_211_19 a_291_70 VDD pmos_3p3 w=34 l=6
X22 a_82_14 a_139_41 a_128_19 GND nmos_3p3 w=17 l=6
X23 a_139_41 CLK GND GND nmos_3p3 w=17 l=6
X24 a_211_19 a_139_41 a_200_70 VDD pmos_3p3 w=34 l=6
X25 a_82_14 CLK a_128_70 VDD pmos_3p3 w=34 l=6
X26 a_139_41 CLK VDD VDD pmos_3p3 w=34 l=6
X27 a_77_19 SN a_41_70 GND nmos_3p3 w=17 l=6
X28 Q QN GND GND nmos_3p3 w=17 l=6
X29 a_234_19 a_139_41 a_211_19 GND nmos_3p3 w=17 l=6
X30 a_172_19 CLK a_82_14 GND nmos_3p3 w=17 l=6
X31 Q QN VDD VDD pmos_3p3 w=34 l=6
X32 GND a_82_14 a_77_19 GND nmos_3p3 w=17 l=6
X33 a_57_70 a_82_14 VDD VDD pmos_3p3 w=34 l=6
X34 a_234_70 CLK a_211_19 VDD pmos_3p3 w=34 l=6
X35 GND a_25_19 a_247_47 GND nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
