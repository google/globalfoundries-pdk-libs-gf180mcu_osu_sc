magic
tech gf180mcuC
timestamp 1661875526
<< nwell >>
rect 0 61 134 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 52 19 58 36
rect 75 19 81 36
rect 91 19 97 36
rect 108 19 114 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 52 70 58 104
rect 75 70 81 104
rect 91 70 97 104
rect 108 70 114 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 19 52 36
rect 58 26 75 36
rect 58 21 64 26
rect 69 21 75 26
rect 58 19 75 21
rect 81 19 91 36
rect 97 33 108 36
rect 97 21 100 33
rect 105 21 108 33
rect 97 19 108 21
rect 114 34 124 36
rect 114 21 117 34
rect 122 21 124 34
rect 114 19 124 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 36 104
rect 25 78 28 102
rect 33 78 36 102
rect 25 70 36 78
rect 42 70 52 104
rect 58 102 75 104
rect 58 97 64 102
rect 69 97 75 102
rect 58 70 75 97
rect 81 70 91 104
rect 97 102 108 104
rect 97 78 100 102
rect 105 78 108 102
rect 97 70 108 78
rect 114 102 124 104
rect 114 72 117 102
rect 122 72 124 102
rect 114 70 124 72
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 64 21 69 26
rect 100 21 105 33
rect 117 21 122 34
<< pdiffc >>
rect 11 72 16 102
rect 28 78 33 102
rect 64 97 69 102
rect 100 78 105 102
rect 117 72 122 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
rect 81 118 90 120
rect 81 113 83 118
rect 88 113 90 118
rect 81 111 90 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
rect 107 113 112 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 52 104 58 109
rect 75 104 81 109
rect 91 104 97 109
rect 108 104 114 109
rect 19 68 25 70
rect 36 68 42 70
rect 19 63 42 68
rect 52 68 58 70
rect 75 68 81 70
rect 52 66 62 68
rect 19 52 25 63
rect 52 61 54 66
rect 60 61 62 66
rect 52 59 62 61
rect 71 66 81 68
rect 71 60 73 66
rect 79 60 81 66
rect 91 68 97 70
rect 108 68 114 70
rect 91 63 114 68
rect 71 58 81 60
rect 19 50 32 52
rect 19 44 24 50
rect 30 44 32 50
rect 19 42 32 44
rect 47 46 58 48
rect 19 38 42 42
rect 47 40 49 46
rect 55 40 58 46
rect 47 38 58 40
rect 19 36 25 38
rect 36 36 42 38
rect 52 36 58 38
rect 75 36 81 58
rect 87 56 97 58
rect 87 51 89 56
rect 95 51 97 56
rect 108 52 114 63
rect 87 49 97 51
rect 91 36 97 49
rect 102 50 114 52
rect 102 44 104 50
rect 110 44 114 50
rect 102 42 114 44
rect 108 36 114 42
rect 19 14 25 19
rect 36 14 42 19
rect 52 14 58 19
rect 75 14 81 19
rect 91 14 97 19
rect 108 14 114 19
<< polycontact >>
rect 54 61 60 66
rect 73 60 79 66
rect 24 44 30 50
rect 49 40 55 46
rect 89 51 95 56
rect 104 44 110 50
<< metal1 >>
rect 0 118 134 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 134 118
rect 0 111 134 112
rect 11 102 16 104
rect 28 102 33 111
rect 64 102 69 104
rect 64 91 69 97
rect 63 89 69 91
rect 100 102 105 111
rect 61 83 63 89
rect 69 83 71 89
rect 28 76 33 78
rect 11 65 16 72
rect 54 73 94 78
rect 100 76 105 78
rect 117 102 122 104
rect 54 66 60 73
rect 89 68 94 73
rect 117 68 122 72
rect 73 66 79 68
rect 11 60 47 65
rect 52 61 54 66
rect 60 61 62 66
rect 11 34 16 60
rect 41 56 47 60
rect 73 56 79 60
rect 89 62 122 68
rect 89 57 95 62
rect 41 51 79 56
rect 87 56 97 57
rect 87 51 89 56
rect 95 51 97 56
rect 22 44 24 50
rect 30 44 32 50
rect 102 46 104 50
rect 47 40 49 46
rect 55 44 104 46
rect 110 44 112 50
rect 55 40 109 44
rect 11 19 16 21
rect 28 34 33 36
rect 63 34 69 35
rect 61 28 63 34
rect 69 28 71 34
rect 100 33 105 35
rect 63 26 69 28
rect 28 12 33 21
rect 64 19 69 21
rect 100 12 105 21
rect 117 34 122 62
rect 117 19 122 21
rect 0 11 134 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 134 11
rect 0 0 134 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 63 83 69 89
rect 24 44 30 50
rect 104 44 110 50
rect 63 28 69 34
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 63 90 69 91
rect 62 89 70 90
rect 62 83 63 89
rect 69 83 70 89
rect 62 82 70 83
rect 23 50 31 51
rect 22 44 24 50
rect 30 44 32 50
rect 23 43 31 44
rect 63 35 69 82
rect 103 50 111 51
rect 102 44 104 50
rect 110 44 112 50
rect 103 43 111 44
rect 61 34 71 35
rect 61 28 63 34
rect 69 28 71 34
rect 61 27 71 28
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 66 85 66 85 1 Y
port 3 n
rlabel metal2 27 47 27 47 1 A
port 1 n
rlabel metal2 107 47 107 47 1 B
port 4 n
<< end >>
