* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_dffsrn_1 D SN RN Q QN CLKN
X0 a_156_109 a_133_14 a_82_14 VDD pmos_3p3 w=34 l=6
X1 VSS a_41_109 a_156_19 VSS nmos_3p3 w=17 l=6
X2 a_82_14 CLKN a_123_109 VDD pmos_3p3 w=34 l=6
X3 a_212_109 CLKN a_195_19 VDD pmos_3p3 w=34 l=6
X4 VSS a_25_19 a_216_68 VSS nmos_3p3 w=17 l=6
X5 a_195_19 CLKN a_184_19 VSS nmos_3p3 w=17 l=6
X6 a_133_14 CLKN VSS VSS nmos_3p3 w=17 l=6
X7 a_216_68 SN a_275_19 VSS nmos_3p3 w=17 l=6
X8 a_25_19 RN VDD VDD pmos_3p3 w=34 l=6
X9 a_123_109 D VDD VDD pmos_3p3 w=34 l=6
X10 VDD a_216_68 QN VDD pmos_3p3 w=34 l=6
X11 Q QN VDD VDD pmos_3p3 w=34 l=6
X12 a_41_109 a_25_19 VSS VSS nmos_3p3 w=17 l=6
X13 a_25_19 RN VSS VSS nmos_3p3 w=17 l=6
X14 a_82_14 a_133_14 a_123_19 VSS nmos_3p3 w=17 l=6
X15 a_256_109 SN VDD VDD pmos_3p3 w=34 l=6
X16 a_275_19 a_195_19 VSS VSS nmos_3p3 w=17 l=6
X17 VDD a_195_19 a_256_109 VDD pmos_3p3 w=34 l=6
X18 a_212_19 a_133_14 a_195_19 VSS nmos_3p3 w=17 l=6
X19 a_216_68 a_25_19 a_256_109 VDD pmos_3p3 w=34 l=6
X20 VSS a_216_68 a_212_19 VSS nmos_3p3 w=17 l=6
X21 a_77_19 SN a_41_109 VSS nmos_3p3 w=17 l=6
X22 a_57_109 a_82_14 VDD VDD pmos_3p3 w=34 l=6
X23 a_57_109 a_25_19 a_41_109 VDD pmos_3p3 w=34 l=6
X24 VDD SN a_57_109 VDD pmos_3p3 w=34 l=6
X25 a_195_19 a_133_14 a_184_109 VDD pmos_3p3 w=34 l=6
X26 Q QN VSS VSS nmos_3p3 w=17 l=6
X27 a_184_109 a_41_109 VDD VDD pmos_3p3 w=34 l=6
X28 VSS a_82_14 a_77_19 VSS nmos_3p3 w=17 l=6
X29 a_156_19 CLKN a_82_14 VSS nmos_3p3 w=17 l=6
X30 VDD a_41_109 a_156_109 VDD pmos_3p3 w=34 l=6
X31 a_133_14 CLKN VDD VDD pmos_3p3 w=34 l=6
X32 a_123_19 D VSS VSS nmos_3p3 w=17 l=6
X33 VDD a_216_68 a_212_109 VDD pmos_3p3 w=34 l=6
X34 a_184_19 a_41_109 VSS VSS nmos_3p3 w=17 l=6
X35 VSS a_216_68 QN VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
