# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_1 0 0 ;
  SIZE 5.35 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 5.35 6.35 ;
        RECT 3.65 3.6 3.9 6.35 ;
        RECT 1.4 4 1.75 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.35 0.7 ;
        RECT 3.65 0 3.9 1.9 ;
        RECT 1.4 0 1.75 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.95 2.95 1.45 3.25 ;
      LAYER Metal2 ;
        RECT 0.95 2.95 1.45 3.25 ;
        RECT 1 2.9 1.4 3.3 ;
      LAYER Via1 ;
        RECT 1.07 2.97 1.33 3.23 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.75 2.3 4.25 2.6 ;
      LAYER Metal2 ;
        RECT 3.75 2.25 4.25 2.65 ;
      LAYER Via1 ;
        RECT 3.87 2.32 4.13 2.58 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 4.15 3.2 4.65 ;
        RECT 2.9 3.5 3.15 5.3 ;
        RECT 2.45 1.65 3.15 1.9 ;
        RECT 2.9 1.05 3.15 1.9 ;
        RECT 2.45 3.5 3.15 3.75 ;
        RECT 2.45 1.65 2.7 3.75 ;
      LAYER Metal2 ;
        RECT 2.8 4.2 3.3 4.6 ;
      LAYER Via1 ;
        RECT 2.92 4.27 3.18 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 3.05 2.9 3.55 3.3 ;
    LAYER Via1 ;
      RECT 3.17 2.97 3.43 3.23 ;
    LAYER Metal1 ;
      RECT 4.5 1.05 4.75 5.3 ;
      RECT 3.05 2.95 4.75 3.25 ;
      RECT 0.55 3.5 0.8 5.3 ;
      RECT 0.45 1.6 0.7 3.9 ;
      RECT 0.45 2.2 2.15 2.5 ;
      RECT 0.55 1.05 0.8 1.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_1
