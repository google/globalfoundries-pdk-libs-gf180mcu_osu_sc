* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsr_1 D Q QN RN SN CLK VDD VSS
X0 a_82_16# CLK a_123_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_212_111# CLK a_195_21# VDD pfet_03p3 w=1.7u l=0.3u
X2 VSS a_41_111# a_156_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_195_21# CLK a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X4 VSS a_25_21# a_216_70# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_133_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
X6 a_216_70# SN a_275_21# VSS nfet_03p3 w=0.85u l=0.3u
X7 a_123_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X8 VDD a_216_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X9 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X10 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X11 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X12 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X13 a_82_16# a_133_16# a_123_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 a_256_111# SN VDD VDD pfet_03p3 w=1.7u l=0.3u
X15 a_275_21# a_195_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X16 VDD a_195_21# a_256_111# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_212_21# a_133_16# a_195_21# VSS nfet_03p3 w=0.85u l=0.3u
X18 a_216_70# a_25_21# a_256_111# VDD pfet_03p3 w=1.7u l=0.3u
X19 VSS a_216_70# a_212_21# VSS nfet_03p3 w=0.85u l=0.3u
X20 a_77_21# SN a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_57_111# a_82_16# VDD VDD pfet_03p3 w=1.7u l=0.3u
X22 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 VDD SN a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X24 a_195_21# a_133_16# a_184_111# VDD pfet_03p3 w=1.7u l=0.3u
X25 VSS a_82_16# a_77_21# VSS nfet_03p3 w=0.85u l=0.3u
X26 a_156_21# CLK a_82_16# VSS nfet_03p3 w=0.85u l=0.3u
X27 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X28 VDD a_41_111# a_156_111# VDD pfet_03p3 w=1.7u l=0.3u
X29 a_184_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X30 a_133_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 a_123_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X32 a_184_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X33 VSS a_216_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X34 a_156_111# a_133_16# a_82_16# VDD pfet_03p3 w=1.7u l=0.3u
X35 VDD a_216_70# a_212_111# VDD pfet_03p3 w=1.7u l=0.3u
.ends
