
.inc "../../char/techfiles/design.hspice"
.lib "../../char/techfiles/sm141064.hspice" typical

.GLOBAL VDD
.GLOBAL GND

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_2
.ends

** hspice subcircuit dictionary
