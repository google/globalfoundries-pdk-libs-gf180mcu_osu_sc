# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tbuf_1 0 0 ;
  SIZE 5.35 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 5.35 6.15 ;
        RECT 3.65 3.5 3.9 6.15 ;
        RECT 1.4 3.9 1.75 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.35 0.6 ;
        RECT 3.65 0 3.9 1.8 ;
        RECT 1.4 0 1.75 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 2.85 1.45 3.15 ;
      LAYER MET2 ;
        RECT 0.95 2.85 1.45 3.15 ;
        RECT 1 2.8 1.4 3.2 ;
      LAYER VIA12 ;
        RECT 1.07 2.87 1.33 3.13 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.75 2.2 4.25 2.5 ;
      LAYER MET2 ;
        RECT 3.75 2.15 4.25 2.55 ;
      LAYER VIA12 ;
        RECT 3.87 2.22 4.13 2.48 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 4.05 3.2 4.55 ;
        RECT 2.9 3.4 3.15 5.2 ;
        RECT 2.45 1.55 3.15 1.8 ;
        RECT 2.9 0.95 3.15 1.8 ;
        RECT 2.45 3.4 3.15 3.65 ;
        RECT 2.45 1.55 2.7 3.65 ;
      LAYER MET2 ;
        RECT 2.8 4.1 3.3 4.5 ;
      LAYER VIA12 ;
        RECT 2.92 4.17 3.18 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 3.05 2.8 3.55 3.2 ;
    LAYER VIA12 ;
      RECT 3.17 2.87 3.43 3.13 ;
    LAYER MET1 ;
      RECT 4.5 0.95 4.75 5.2 ;
      RECT 3.05 2.85 4.75 3.15 ;
      RECT 0.55 3.4 0.8 5.2 ;
      RECT 0.45 1.5 0.7 3.8 ;
      RECT 0.45 2.1 2.15 2.4 ;
      RECT 0.55 0.95 0.8 1.8 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tbuf_1
