VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_addh_1 0 0 ;
  SIZE 8.6 BY 6.15 ;
  SYMMETRY X Y ;
  SITE 9T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 2.2 4.4 2.5 ;
        RECT 1.5 2.2 2 2.5 ;
      LAYER MET2 ;
        RECT 3.9 2.15 4.4 2.55 ;
        RECT 1.5 2.2 4.4 2.5 ;
        RECT 1.5 2.15 2 2.55 ;
      LAYER VIA12 ;
        RECT 1.62 2.22 1.88 2.48 ;
        RECT 4.02 2.22 4.28 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 1.9 5.5 2.4 ;
        RECT 2.35 2.15 2.85 2.45 ;
        RECT 2.35 1.55 2.85 1.85 ;
        RECT 2.45 1.55 2.75 2.45 ;
      LAYER MET2 ;
        RECT 5.15 1.95 5.55 2.35 ;
        RECT 5.2 1.55 5.5 2.4 ;
        RECT 5.15 1.55 5.5 2.35 ;
        RECT 2.35 1.55 5.5 1.85 ;
        RECT 2.4 1.5 2.8 1.9 ;
      LAYER VIA12 ;
        RECT 2.47 1.57 2.73 1.83 ;
        RECT 5.22 2.02 5.48 2.28 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
        RECT 0.55 0.95 0.8 5.2 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END CO
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.6 0.6 ;
        RECT 6.65 0 6.9 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
      LAYER MET2 ;
        RECT 6.7 0.25 7.2 0.55 ;
        RECT 6.75 0.2 7.15 0.6 ;
        RECT 5.25 0.25 5.75 0.55 ;
        RECT 5.3 0.2 5.7 0.6 ;
        RECT 4.05 0.25 4.55 0.55 ;
        RECT 4.1 0.2 4.5 0.6 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
        RECT 4.17 0.27 4.43 0.53 ;
        RECT 5.37 0.27 5.63 0.53 ;
        RECT 6.82 0.27 7.08 0.53 ;
    END
  END GND
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.7 2.85 8.2 3.15 ;
        RECT 7.75 2.8 8.1 3.2 ;
        RECT 7.5 3.5 8 5.2 ;
        RECT 7.75 0.95 8 5.2 ;
      LAYER MET2 ;
        RECT 7.7 2.8 8.2 3.2 ;
      LAYER VIA12 ;
        RECT 7.82 2.87 8.08 3.13 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.6 6.15 ;
        RECT 6.65 4.5 6.9 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
      LAYER MET2 ;
        RECT 6.45 5.6 6.95 5.9 ;
        RECT 6.5 5.55 6.9 5.95 ;
        RECT 5.25 5.6 5.75 5.9 ;
        RECT 5.3 5.55 5.7 5.95 ;
        RECT 4.05 5.6 4.55 5.9 ;
        RECT 4.1 5.55 4.5 5.95 ;
        RECT 2.85 5.6 3.35 5.9 ;
        RECT 2.9 5.55 3.3 5.95 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
        RECT 2.97 5.62 3.23 5.88 ;
        RECT 4.17 5.62 4.43 5.88 ;
        RECT 5.37 5.62 5.63 5.88 ;
        RECT 6.57 5.62 6.83 5.88 ;
    END
  END VDD
  OBS
    LAYER MET2 ;
      RECT 6.3 2.95 6.8 3.35 ;
      RECT 3 2.9 3.5 3.3 ;
      RECT 3 2.95 6.8 3.25 ;
    LAYER VIA12 ;
      RECT 6.42 3.02 6.68 3.28 ;
      RECT 3.12 2.97 3.38 3.23 ;
    LAYER MET1 ;
      RECT 5.55 3.5 6.05 5.2 ;
      RECT 5.55 2.75 5.8 5.2 ;
      RECT 4.7 2.75 6.05 3 ;
      RECT 5.75 2.5 6.75 2.75 ;
      RECT 4.7 1.35 4.95 3 ;
      RECT 6.5 2.2 7.25 2.5 ;
      RECT 5.55 0.85 5.8 1.45 ;
      RECT 3.85 0.85 4.1 1.45 ;
      RECT 3.85 0.85 5.8 1.1 ;
      RECT 2.25 2.95 2.5 5.2 ;
      RECT 1.05 2.95 3.5 3.25 ;
      RECT 3.1 0.95 3.35 3.25 ;
      RECT 6.3 3 6.8 3.3 ;
  END
END gf180mcu_osu_sc_9T_addh_1
