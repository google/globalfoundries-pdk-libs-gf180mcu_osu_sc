# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_and2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_and2_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 2.25 5.45 2.5 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 2.1 0 2.5 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 2.85 2.4 3.15 ;
      LAYER MET2 ;
        RECT 1.9 2.8 2.4 3.2 ;
      LAYER VIA12 ;
        RECT 2.02 2.87 2.28 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 4.85 3.6 5.15 ;
        RECT 3.1 4.8 3.5 5.15 ;
        RECT 3.1 4.8 3.45 5.2 ;
        RECT 3.1 0.95 3.35 7.15 ;
      LAYER MET2 ;
        RECT 3.1 4.8 3.6 5.2 ;
      LAYER VIA12 ;
        RECT 3.22 4.87 3.48 5.13 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.35 4.1 2.85 4.5 ;
      RECT 1.3 4.1 1.8 4.5 ;
    LAYER VIA12 ;
      RECT 2.47 4.17 2.73 4.43 ;
      RECT 1.42 4.17 1.68 4.43 ;
    LAYER MET1 ;
      RECT 1.4 1.9 1.65 7.15 ;
      RECT 1.3 4.15 2.85 4.45 ;
      RECT 0.7 1.9 1.65 2.15 ;
      RECT 0.7 0.95 0.95 2.15 ;
  END
END gf180mcu_osu_sc_12T_and2_1
