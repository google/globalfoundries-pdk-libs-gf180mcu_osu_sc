# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tieh
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tieh 0 0 ;
  SIZE 2.2 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 2.2 6.35 ;
        RECT 0.55 3.6 0.8 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 2.2 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.3 3.6 1.8 3.9 ;
        RECT 1.4 3.55 1.65 5.3 ;
      LAYER Metal2 ;
        RECT 1.3 3.55 1.8 3.95 ;
      LAYER Via1 ;
        RECT 1.42 3.62 1.68 3.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.15 2.3 1.65 2.55 ;
      RECT 1.4 1.05 1.65 2.55 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tieh
