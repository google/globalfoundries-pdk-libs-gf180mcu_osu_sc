# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__antfill
  CLASS CORE ;
  ORIGIN 0 0.05 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__antfill 0 -0.05 ;
  SIZE 2.2 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.6 2.2 6.3 ;
        RECT 1.4 3.55 1.65 6.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.05 2.2 0.65 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 2.25 1.65 2.55 ;
        RECT 1.4 1 1.65 2.55 ;
        RECT 0.55 1 0.8 5.25 ;
        RECT 0.5 2.2 0.8 2.65 ;
      LAYER Metal2 ;
        RECT 0.45 2.25 0.95 2.55 ;
        RECT 0.5 2.2 0.9 2.6 ;
      LAYER Via1 ;
        RECT 0.57 2.27 0.83 2.53 ;
    END
  END A
END gf180mcu_osu_sc_gp9t3v3__antfill
