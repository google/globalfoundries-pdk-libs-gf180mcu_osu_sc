magic
tech gf180mcuC
timestamp 1661874254
<< nwell >>
rect 0 61 280 123
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 53 19 59 36
rect 70 19 76 36
rect 87 19 93 36
rect 104 19 110 36
rect 121 19 127 36
rect 138 19 144 36
rect 155 19 161 36
rect 172 19 178 36
rect 189 19 195 36
rect 206 19 212 36
rect 223 19 229 36
rect 255 19 261 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 53 70 59 104
rect 70 70 76 104
rect 87 70 93 104
rect 104 70 110 104
rect 121 70 127 104
rect 138 70 144 104
rect 155 70 161 104
rect 172 70 178 104
rect 189 70 195 104
rect 206 70 212 104
rect 223 70 229 104
rect 255 70 261 104
<< ndiff >>
rect 9 26 19 36
rect 9 21 11 26
rect 16 21 19 26
rect 9 19 19 21
rect 25 26 36 36
rect 25 21 28 26
rect 33 21 36 26
rect 25 19 36 21
rect 42 26 53 36
rect 42 21 45 26
rect 50 21 53 26
rect 42 19 53 21
rect 59 26 70 36
rect 59 21 62 26
rect 67 21 70 26
rect 59 19 70 21
rect 76 19 87 36
rect 93 26 104 36
rect 93 21 96 26
rect 101 21 104 26
rect 93 19 104 21
rect 110 26 121 36
rect 110 21 113 26
rect 118 21 121 26
rect 110 19 121 21
rect 127 26 138 36
rect 127 21 130 26
rect 135 21 138 26
rect 127 19 138 21
rect 144 26 155 36
rect 144 21 147 26
rect 152 21 155 26
rect 144 19 155 21
rect 161 26 172 36
rect 161 21 164 26
rect 169 21 172 26
rect 161 19 172 21
rect 178 19 189 36
rect 195 19 206 36
rect 212 26 223 36
rect 212 21 215 26
rect 220 21 223 26
rect 212 19 223 21
rect 229 26 239 36
rect 229 21 232 26
rect 237 21 239 26
rect 229 19 239 21
rect 245 26 255 36
rect 245 21 247 26
rect 252 21 255 26
rect 245 19 255 21
rect 261 26 271 36
rect 261 21 264 26
rect 269 21 271 26
rect 261 19 271 21
<< pdiff >>
rect 9 102 19 104
rect 9 96 11 102
rect 16 96 19 102
rect 9 70 19 96
rect 25 102 36 104
rect 25 96 28 102
rect 33 96 36 102
rect 25 70 36 96
rect 42 102 53 104
rect 42 96 45 102
rect 50 96 53 102
rect 42 70 53 96
rect 59 102 70 104
rect 59 97 62 102
rect 67 97 70 102
rect 59 70 70 97
rect 76 70 87 104
rect 93 102 104 104
rect 93 96 96 102
rect 101 96 104 102
rect 93 70 104 96
rect 110 102 121 104
rect 110 96 113 102
rect 118 96 121 102
rect 110 70 121 96
rect 127 102 138 104
rect 127 96 130 102
rect 135 96 138 102
rect 127 70 138 96
rect 144 102 155 104
rect 144 96 147 102
rect 152 96 155 102
rect 144 70 155 96
rect 161 89 172 104
rect 161 83 164 89
rect 169 83 172 89
rect 161 70 172 83
rect 178 70 189 104
rect 195 70 206 104
rect 212 102 223 104
rect 212 96 215 102
rect 220 96 223 102
rect 212 70 223 96
rect 229 102 239 104
rect 229 96 232 102
rect 237 96 239 102
rect 229 70 239 96
rect 245 102 255 104
rect 245 96 247 102
rect 252 96 255 102
rect 245 70 255 96
rect 261 102 271 104
rect 261 96 264 102
rect 269 96 271 102
rect 261 70 271 96
<< ndiffc >>
rect 11 21 16 26
rect 28 21 33 26
rect 45 21 50 26
rect 62 21 67 26
rect 96 21 101 26
rect 113 21 118 26
rect 130 21 135 26
rect 147 21 152 26
rect 164 21 169 26
rect 215 21 220 26
rect 232 21 237 26
rect 247 21 252 26
rect 264 21 269 26
<< pdiffc >>
rect 11 96 16 102
rect 28 96 33 102
rect 45 96 50 102
rect 62 97 67 102
rect 96 96 101 102
rect 113 96 118 102
rect 130 96 135 102
rect 147 96 152 102
rect 164 83 169 89
rect 215 96 220 102
rect 232 96 237 102
rect 247 96 252 102
rect 264 96 269 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 129 10 138 12
rect 129 5 131 10
rect 136 5 138 10
rect 129 3 138 5
rect 153 10 162 12
rect 153 5 155 10
rect 160 5 162 10
rect 153 3 162 5
rect 177 10 186 12
rect 177 5 179 10
rect 184 5 186 10
rect 177 3 186 5
rect 201 10 210 12
rect 201 5 203 10
rect 208 5 210 10
rect 201 3 210 5
rect 225 10 234 12
rect 225 5 227 10
rect 232 5 234 10
rect 225 3 234 5
rect 249 10 258 12
rect 249 5 251 10
rect 256 5 258 10
rect 249 3 258 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
rect 81 118 90 120
rect 81 113 83 118
rect 88 113 90 118
rect 81 111 90 113
rect 105 118 114 120
rect 105 113 107 118
rect 112 113 114 118
rect 105 111 114 113
rect 129 118 138 120
rect 129 113 131 118
rect 136 113 138 118
rect 129 111 138 113
rect 153 118 162 120
rect 153 113 155 118
rect 160 113 162 118
rect 153 111 162 113
rect 177 118 186 120
rect 177 113 179 118
rect 184 113 186 118
rect 177 111 186 113
rect 201 118 210 120
rect 201 113 203 118
rect 208 113 210 118
rect 201 111 210 113
rect 225 118 234 120
rect 225 113 227 118
rect 232 113 234 118
rect 225 111 234 113
rect 249 118 258 120
rect 249 113 251 118
rect 256 113 258 118
rect 249 111 258 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
rect 131 5 136 10
rect 155 5 160 10
rect 179 5 184 10
rect 203 5 208 10
rect 227 5 232 10
rect 251 5 256 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
rect 83 113 88 118
rect 107 113 112 118
rect 131 113 136 118
rect 155 113 160 118
rect 179 113 184 118
rect 203 113 208 118
rect 227 113 232 118
rect 251 113 256 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 53 104 59 109
rect 70 104 76 109
rect 87 104 93 109
rect 104 104 110 109
rect 121 104 127 109
rect 138 104 144 109
rect 155 104 161 109
rect 172 104 178 109
rect 189 104 195 109
rect 206 104 212 109
rect 223 104 229 109
rect 255 104 261 109
rect 19 52 25 70
rect 36 65 42 70
rect 30 63 42 65
rect 30 57 32 63
rect 38 57 42 63
rect 30 55 42 57
rect 12 50 25 52
rect 12 44 14 50
rect 20 44 25 50
rect 12 42 25 44
rect 19 36 25 42
rect 36 36 42 55
rect 53 52 59 70
rect 70 68 76 70
rect 87 68 93 70
rect 104 68 110 70
rect 121 68 127 70
rect 70 66 82 68
rect 70 60 74 66
rect 80 60 82 66
rect 70 58 82 60
rect 87 63 110 68
rect 115 66 127 68
rect 51 50 61 52
rect 51 44 53 50
rect 59 44 61 50
rect 51 42 61 44
rect 53 36 59 42
rect 70 36 76 58
rect 87 55 93 63
rect 115 60 117 66
rect 123 60 127 66
rect 115 58 127 60
rect 87 53 102 55
rect 87 47 94 53
rect 100 47 102 53
rect 87 45 102 47
rect 87 40 110 45
rect 87 36 93 40
rect 104 36 110 40
rect 121 36 127 58
rect 138 55 144 70
rect 155 55 161 70
rect 172 55 178 70
rect 189 68 195 70
rect 189 66 201 68
rect 189 60 193 66
rect 199 60 201 66
rect 189 58 201 60
rect 138 53 149 55
rect 138 47 141 53
rect 147 47 149 53
rect 138 45 149 47
rect 155 53 166 55
rect 155 47 158 53
rect 164 47 166 53
rect 155 45 166 47
rect 172 53 184 55
rect 172 47 176 53
rect 182 47 184 53
rect 172 45 184 47
rect 138 36 144 45
rect 155 36 161 45
rect 172 36 178 45
rect 189 36 195 58
rect 206 53 212 70
rect 223 55 229 70
rect 255 55 261 70
rect 202 51 212 53
rect 202 45 204 51
rect 210 45 212 51
rect 217 53 229 55
rect 217 47 219 53
rect 225 47 229 53
rect 217 45 229 47
rect 249 53 261 55
rect 249 47 251 53
rect 257 47 261 53
rect 249 45 261 47
rect 202 43 212 45
rect 206 36 212 43
rect 223 36 229 45
rect 255 36 261 45
rect 19 14 25 19
rect 36 14 42 19
rect 53 14 59 19
rect 70 14 76 19
rect 87 14 93 19
rect 104 14 110 19
rect 121 14 127 19
rect 138 14 144 19
rect 155 14 161 19
rect 172 14 178 19
rect 189 14 195 19
rect 206 14 212 19
rect 223 14 229 19
rect 255 14 261 19
<< polycontact >>
rect 32 57 38 63
rect 14 44 20 50
rect 74 60 80 66
rect 53 44 59 50
rect 117 60 123 66
rect 94 47 100 53
rect 193 60 199 66
rect 141 47 147 53
rect 158 47 164 53
rect 176 47 182 53
rect 204 45 210 51
rect 219 47 225 53
rect 251 47 257 53
<< metal1 >>
rect 0 118 280 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 83 118
rect 89 112 107 118
rect 113 112 131 118
rect 137 112 155 118
rect 161 112 179 118
rect 185 112 203 118
rect 209 112 227 118
rect 233 112 251 118
rect 257 112 280 118
rect 0 111 280 112
rect 11 102 16 104
rect 11 89 16 96
rect 28 102 33 111
rect 28 94 33 96
rect 45 102 50 104
rect 45 89 50 96
rect 62 102 68 104
rect 62 94 68 96
rect 96 102 101 111
rect 96 94 101 96
rect 113 102 118 104
rect 11 84 50 89
rect 113 89 118 96
rect 130 102 135 111
rect 130 94 135 96
rect 147 102 152 104
rect 147 89 152 96
rect 215 102 220 111
rect 215 94 220 96
rect 232 102 237 104
rect 113 84 152 89
rect 162 83 164 89
rect 170 83 172 89
rect 32 73 80 79
rect 32 63 38 73
rect 32 55 38 57
rect 43 62 69 68
rect 43 50 48 62
rect 64 53 69 62
rect 74 66 80 73
rect 117 72 199 78
rect 117 66 123 72
rect 80 60 117 66
rect 74 58 80 60
rect 117 58 123 60
rect 128 61 182 67
rect 128 53 134 61
rect 12 44 14 50
rect 20 44 48 50
rect 53 50 59 52
rect 64 47 94 53
rect 100 47 134 53
rect 141 53 147 55
rect 176 53 182 61
rect 193 66 199 72
rect 193 58 199 60
rect 232 67 237 96
rect 247 102 252 111
rect 247 94 252 96
rect 264 102 269 104
rect 264 67 269 96
rect 232 66 238 67
rect 264 66 273 67
rect 232 60 233 66
rect 239 60 241 66
rect 264 60 267 66
rect 273 60 275 66
rect 232 59 238 60
rect 264 59 273 60
rect 156 47 158 53
rect 164 47 166 53
rect 174 47 176 53
rect 182 47 184 53
rect 53 42 59 44
rect 141 42 147 47
rect 195 45 204 51
rect 210 45 212 51
rect 217 47 219 53
rect 225 47 227 53
rect 195 42 201 45
rect 53 36 201 42
rect 10 27 16 29
rect 10 19 16 21
rect 28 26 33 28
rect 28 12 33 21
rect 44 27 50 29
rect 44 19 50 21
rect 62 27 68 29
rect 62 19 68 21
rect 96 26 101 28
rect 96 12 101 21
rect 113 27 119 29
rect 113 19 119 21
rect 130 26 135 28
rect 130 12 135 21
rect 146 27 152 29
rect 146 19 152 21
rect 164 27 170 29
rect 164 19 170 21
rect 215 26 220 28
rect 215 12 220 21
rect 232 26 237 59
rect 249 47 251 53
rect 257 47 259 53
rect 232 19 237 21
rect 247 26 252 28
rect 247 12 252 21
rect 264 26 269 59
rect 264 19 269 21
rect 0 11 280 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 131 11
rect 137 5 155 11
rect 161 5 179 11
rect 185 5 203 11
rect 209 5 227 11
rect 233 5 251 11
rect 257 5 280 11
rect 0 0 280 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 83 113 88 118
rect 88 113 89 118
rect 83 112 89 113
rect 107 113 112 118
rect 112 113 113 118
rect 107 112 113 113
rect 131 113 136 118
rect 136 113 137 118
rect 131 112 137 113
rect 155 113 160 118
rect 160 113 161 118
rect 155 112 161 113
rect 179 113 184 118
rect 184 113 185 118
rect 179 112 185 113
rect 203 113 208 118
rect 208 113 209 118
rect 203 112 209 113
rect 227 113 232 118
rect 232 113 233 118
rect 227 112 233 113
rect 251 113 256 118
rect 256 113 257 118
rect 251 112 257 113
rect 62 97 67 102
rect 67 97 68 102
rect 62 96 68 97
rect 164 83 169 89
rect 169 83 170 89
rect 32 57 38 63
rect 14 44 20 50
rect 53 44 59 50
rect 233 60 239 66
rect 267 60 273 66
rect 158 47 164 53
rect 219 47 225 53
rect 10 26 16 27
rect 10 21 11 26
rect 11 21 16 26
rect 44 26 50 27
rect 44 21 45 26
rect 45 21 50 26
rect 62 26 68 27
rect 62 21 67 26
rect 67 21 68 26
rect 113 26 119 27
rect 113 21 118 26
rect 118 21 119 26
rect 146 26 152 27
rect 146 21 147 26
rect 147 21 152 26
rect 164 26 170 27
rect 164 21 169 26
rect 169 21 170 26
rect 251 47 257 53
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 131 10 137 11
rect 131 5 136 10
rect 136 5 137 10
rect 155 10 161 11
rect 155 5 160 10
rect 160 5 161 10
rect 179 10 185 11
rect 179 5 184 10
rect 184 5 185 10
rect 203 10 209 11
rect 203 5 208 10
rect 208 5 209 10
rect 227 10 233 11
rect 227 5 232 10
rect 232 5 233 10
rect 251 10 257 11
rect 251 5 256 10
rect 256 5 257 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 81 112 83 118
rect 89 112 91 118
rect 105 112 107 118
rect 113 112 115 118
rect 129 112 131 118
rect 137 112 139 118
rect 153 112 155 118
rect 161 112 163 118
rect 177 112 179 118
rect 185 112 187 118
rect 201 112 203 118
rect 209 112 211 118
rect 225 112 227 118
rect 233 112 235 118
rect 249 112 251 118
rect 257 112 259 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 62 103 68 104
rect 61 102 69 103
rect 60 96 62 102
rect 68 96 257 102
rect 61 95 69 96
rect 31 63 39 64
rect 30 57 32 63
rect 38 57 40 63
rect 31 56 39 57
rect 75 53 81 96
rect 163 89 171 90
rect 162 83 164 89
rect 170 83 225 89
rect 163 82 171 83
rect 157 53 165 54
rect 12 50 22 51
rect 52 50 60 51
rect 12 44 14 50
rect 20 44 22 50
rect 51 44 53 50
rect 59 44 61 50
rect 75 47 158 53
rect 164 47 166 53
rect 12 43 22 44
rect 52 43 60 44
rect 10 28 16 29
rect 44 28 50 29
rect 62 28 68 29
rect 9 27 17 28
rect 43 27 51 28
rect 9 21 10 27
rect 16 21 44 27
rect 50 21 51 27
rect 9 20 17 21
rect 43 20 51 21
rect 61 27 69 28
rect 75 27 81 47
rect 157 46 165 47
rect 113 28 119 29
rect 146 28 152 29
rect 61 21 62 27
rect 68 21 81 27
rect 112 27 120 28
rect 145 27 153 28
rect 163 27 171 28
rect 177 27 183 83
rect 219 54 225 83
rect 232 66 240 67
rect 231 60 233 66
rect 239 60 241 66
rect 232 59 240 60
rect 251 54 257 96
rect 266 66 274 67
rect 265 60 267 66
rect 273 60 275 66
rect 266 59 274 60
rect 218 53 226 54
rect 250 53 258 54
rect 218 47 219 53
rect 225 47 226 53
rect 249 47 251 53
rect 257 47 259 53
rect 218 46 226 47
rect 250 46 258 47
rect 219 45 225 46
rect 251 45 257 46
rect 112 21 113 27
rect 119 21 146 27
rect 152 21 153 27
rect 162 21 164 27
rect 170 21 183 27
rect 61 20 69 21
rect 112 20 120 21
rect 145 20 153 21
rect 163 20 171 21
rect 10 19 16 20
rect 44 19 50 20
rect 62 19 68 20
rect 113 19 119 20
rect 146 19 152 20
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 129 5 131 11
rect 137 5 139 11
rect 153 5 155 11
rect 161 5 163 11
rect 177 5 179 11
rect 185 5 187 11
rect 201 5 203 11
rect 209 5 211 11
rect 225 5 227 11
rect 233 5 235 11
rect 249 5 251 11
rect 257 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 17 47 17 47 1 A
port 7 n
rlabel metal2 35 60 35 60 1 B
port 8 n
rlabel metal2 56 47 56 47 1 CI
port 9 n
rlabel metal2 236 63 236 63 1 S
port 10 n
rlabel metal2 270 63 270 63 1 CO
port 11 n
<< end >>
