VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_tielo
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_tielo 0 0 ;
  SIZE 2.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE 9T ;
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.2 0.6 ;
        RECT 0.55 0 0.8 1.8 ;
      LAYER MET2 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 2.2 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
      LAYER MET2 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 1.55 1.8 1.85 ;
        RECT 1.4 0.95 1.65 1.9 ;
      LAYER MET2 ;
        RECT 1.3 1.5 1.8 1.9 ;
      LAYER VIA12 ;
        RECT 1.42 1.57 1.68 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 2.9 1.65 5.2 ;
      RECT 1.15 2.9 1.65 3.15 ;
  END
END gf180mcu_osu_sc_9T_tielo
