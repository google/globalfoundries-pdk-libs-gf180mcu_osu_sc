# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__addf_1 0 0 ;
  SIZE 14 BY 8.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 14 8.35 ;
        RECT 12.35 5.55 12.6 8.35 ;
        RECT 10.75 5.55 11 8.35 ;
        RECT 6.5 5.55 6.75 8.35 ;
        RECT 4.8 5.55 5.05 8.35 ;
        RECT 1.4 5.55 1.65 8.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14 0.7 ;
        RECT 12.35 0 12.6 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 6.5 0 6.75 1.55 ;
        RECT 4.8 0 5.05 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.7 3.6 9.2 3.9 ;
        RECT 4.6 3.6 5.1 3.9 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.6 9.2 3.9 ;
        RECT 8.75 3.55 9.15 3.95 ;
        RECT 4.65 3.55 5.05 3.95 ;
        RECT 0.65 3.55 1.05 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
        RECT 4.72 3.62 4.98 3.88 ;
        RECT 8.82 3.62 9.08 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.55 4.25 10.05 4.55 ;
        RECT 3.6 4.25 6.25 4.55 ;
        RECT 1.5 4.25 2 4.55 ;
      LAYER Metal2 ;
        RECT 5.75 4.25 10.05 4.55 ;
        RECT 9.6 4.2 10 4.6 ;
        RECT 5.8 4.2 6.2 4.6 ;
        RECT 1.5 4.25 4.1 4.55 ;
        RECT 3.65 4.2 4.05 4.6 ;
        RECT 1.55 4.2 1.95 4.6 ;
      LAYER Via1 ;
        RECT 1.62 4.27 1.88 4.53 ;
        RECT 3.72 4.27 3.98 4.53 ;
        RECT 5.87 4.27 6.13 4.53 ;
        RECT 9.67 4.27 9.93 4.53 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.05 2.3 10.55 2.6 ;
        RECT 6.65 2.3 7.15 2.6 ;
        RECT 2.35 2.95 2.85 3.25 ;
      LAYER Metal2 ;
        RECT 2.45 2.3 10.55 2.6 ;
        RECT 10.1 2.25 10.5 2.65 ;
        RECT 10.15 2.2 10.45 2.65 ;
        RECT 6.7 2.25 7.1 2.65 ;
        RECT 6.75 2.2 7.05 2.65 ;
        RECT 2.35 2.95 2.85 3.25 ;
        RECT 2.4 2.9 2.8 3.3 ;
        RECT 2.45 2.3 2.75 3.3 ;
      LAYER Via1 ;
        RECT 2.47 2.97 2.73 3.23 ;
        RECT 6.77 2.32 7.03 2.58 ;
        RECT 10.17 2.32 10.43 2.58 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.2 2.95 13.75 3.25 ;
        RECT 13.2 2.9 13.6 3.3 ;
        RECT 13.2 1.05 13.45 7.25 ;
      LAYER Metal2 ;
        RECT 13.25 2.95 13.75 3.25 ;
        RECT 13.3 2.9 13.7 3.3 ;
      LAYER Via1 ;
        RECT 13.37 2.97 13.63 3.23 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.6 4.25 12 4.55 ;
        RECT 11.6 1.05 11.85 7.25 ;
      LAYER Metal2 ;
        RECT 11.5 4.25 12 4.55 ;
        RECT 11.55 4.2 11.95 4.6 ;
      LAYER Via1 ;
        RECT 11.62 4.27 11.88 4.53 ;
    END
  END S
  OBS
    LAYER Metal2 ;
      RECT 12.5 2.9 12.9 3.3 ;
      RECT 7.5 2.9 7.9 3.3 ;
      RECT 7.45 2.95 12.95 3.25 ;
      RECT 12.55 2.85 12.85 3.3 ;
    LAYER Via1 ;
      RECT 12.57 2.97 12.83 3.23 ;
      RECT 7.57 2.97 7.83 3.23 ;
    LAYER Metal1 ;
      RECT 8.2 1.05 8.45 7.25 ;
      RECT 8.2 2.95 11.35 3.25 ;
      RECT 3.1 1.05 3.35 7.25 ;
      RECT 3.1 2.95 7.95 3.25 ;
      RECT 5.65 1.8 7.6 2.05 ;
      RECT 7.35 1.05 7.6 2.05 ;
      RECT 5.65 1.05 5.9 2.05 ;
      RECT 7.35 5.05 7.6 7.25 ;
      RECT 5.65 5.05 5.9 7.25 ;
      RECT 5.65 5.05 7.6 5.3 ;
      RECT 0.55 2.15 2.5 2.4 ;
      RECT 2.25 1.05 2.5 2.4 ;
      RECT 0.55 1.05 0.8 2.4 ;
      RECT 2.25 5.05 2.5 7.25 ;
      RECT 0.55 5.05 0.8 7.25 ;
      RECT 0.55 5.05 2.5 5.3 ;
      RECT 12.45 2.95 12.95 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__addf_1
