# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsr_1 0 0 ;
  SIZE 18.7 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 18.7 8.3 ;
        RECT 17.05 5.55 17.3 8.3 ;
        RECT 13.75 6.8 14 8.3 ;
        RECT 11.3 6.3 11.55 8.3 ;
        RECT 8.5 5.55 8.75 8.3 ;
        RECT 5.45 5.55 5.7 8.3 ;
        RECT 3.85 6.3 4.1 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 18.7 0.7 ;
        RECT 17.05 0 17.3 1.9 ;
        RECT 15.3 0 15.55 1.9 ;
        RECT 13.05 0 13.3 1.9 ;
        RECT 11.3 0 11.55 1.9 ;
        RECT 8.5 0 8.75 1.5 ;
        RECT 5.45 0 5.7 1.9 ;
        RECT 4.55 0 4.8 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 11.7 4.25 12.2 4.55 ;
        RECT 9.55 4.25 10.6 4.55 ;
        RECT 9.45 2.25 9.95 2.55 ;
        RECT 9.55 2.25 9.85 4.55 ;
        RECT 6.65 4.25 7.8 4.55 ;
        RECT 7.3 2.3 7.8 2.6 ;
        RECT 7.4 2.3 7.7 4.55 ;
      LAYER Metal2 ;
        RECT 7.3 4.25 12.2 4.55 ;
        RECT 11.75 4.2 12.15 4.6 ;
        RECT 10.1 4.2 10.6 4.6 ;
        RECT 7.3 4.2 7.75 4.6 ;
      LAYER Via1 ;
        RECT 7.42 4.27 7.68 4.53 ;
        RECT 10.22 4.27 10.48 4.53 ;
        RECT 11.82 4.27 12.08 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.95 3.6 6.45 3.9 ;
      LAYER Metal2 ;
        RECT 5.95 3.55 6.45 3.95 ;
      LAYER Via1 ;
        RECT 6.07 3.62 6.33 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17.9 4.9 18.4 5.25 ;
        RECT 17.9 4.85 18.35 5.25 ;
        RECT 17.9 1.05 18.15 7.25 ;
      LAYER Metal2 ;
        RECT 17.9 4.9 18.4 5.2 ;
        RECT 17.95 4.85 18.35 5.25 ;
      LAYER Via1 ;
        RECT 18.02 4.92 18.28 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.2 4.25 17.65 4.55 ;
        RECT 17.3 2.15 17.55 4.55 ;
        RECT 16.2 2.15 17.55 2.4 ;
        RECT 16.2 4.25 16.45 7.25 ;
        RECT 16.2 1.05 16.45 2.4 ;
      LAYER Metal2 ;
        RECT 17.15 4.25 17.65 4.55 ;
        RECT 17.2 4.2 17.6 4.6 ;
      LAYER Via1 ;
        RECT 17.27 4.27 17.53 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.95 4.25 14.45 4.55 ;
        RECT 3.4 4.25 3.9 4.55 ;
      LAYER Metal2 ;
        RECT 13.95 4.2 14.45 4.6 ;
        RECT 3.5 5.55 14.35 5.85 ;
        RECT 14.05 4.2 14.35 5.85 ;
        RECT 3.4 4.2 3.9 4.6 ;
        RECT 3.5 4.2 3.8 5.85 ;
      LAYER Via1 ;
        RECT 3.52 4.27 3.78 4.53 ;
        RECT 14.07 4.27 14.33 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 16.45 2.9 16.85 3.3 ;
      RECT 16.1 2.95 16.9 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 14.85 2.2 15.45 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 14.85 1 15.15 2.6 ;
      RECT 2.75 1 15.15 1.3 ;
      RECT 12.95 2.2 13.45 2.6 ;
      RECT 12.95 1.65 13.35 2.6 ;
      RECT 9.85 1.6 10.25 2 ;
      RECT 9.8 1.65 13.35 1.95 ;
      RECT 13 4.85 13.4 5.25 ;
      RECT 10.8 4.85 11.2 5.25 ;
      RECT 10.75 4.9 13.45 5.2 ;
      RECT 12.1 2.9 12.5 3.3 ;
      RECT 10.15 2.9 10.55 3.3 ;
      RECT 10.1 2.95 12.6 3.25 ;
      RECT 10.85 3.55 11.25 3.95 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 8.15 2.25 8.55 2.65 ;
      RECT 4.4 2.25 4.9 2.65 ;
      RECT 4.4 2.3 8.6 2.6 ;
      RECT 15.35 4.85 15.85 5.25 ;
      RECT 4.4 3.55 4.9 3.95 ;
    LAYER Via1 ;
      RECT 16.52 2.97 16.78 3.23 ;
      RECT 15.47 4.92 15.73 5.18 ;
      RECT 15.07 2.27 15.33 2.53 ;
      RECT 13.07 2.27 13.33 2.53 ;
      RECT 13.07 4.92 13.33 5.18 ;
      RECT 12.17 2.97 12.43 3.23 ;
      RECT 10.92 3.62 11.18 3.88 ;
      RECT 10.87 4.92 11.13 5.18 ;
      RECT 10.22 2.97 10.48 3.23 ;
      RECT 9.92 1.67 10.18 1.93 ;
      RECT 8.22 2.32 8.48 2.58 ;
      RECT 4.52 2.32 4.78 2.58 ;
      RECT 4.52 3.62 4.78 3.88 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 15.45 2.95 15.7 7.25 ;
      RECT 13.05 4.8 13.35 5.3 ;
      RECT 13.05 4.9 15.85 5.2 ;
      RECT 14.45 2.95 16.9 3.25 ;
      RECT 14.45 1.05 14.7 3.25 ;
      RECT 14.6 6.3 14.85 7.25 ;
      RECT 12.9 6.3 13.15 7.25 ;
      RECT 12.9 6.3 14.85 6.55 ;
      RECT 12.15 4.85 12.4 7.25 ;
      RECT 12.15 4.85 12.7 5.1 ;
      RECT 12.45 3.65 12.7 5.1 ;
      RECT 12.15 2.85 12.45 3.9 ;
      RECT 12.15 1.05 12.4 3.9 ;
      RECT 10.75 4.9 11.25 5.2 ;
      RECT 10.85 3.6 11.15 5.2 ;
      RECT 10.8 3.6 11.3 3.9 ;
      RECT 9.9 6.05 10.15 7.25 ;
      RECT 9 6.05 10.15 6.3 ;
      RECT 9 3.55 9.25 6.3 ;
      RECT 8.95 1.7 9.2 3.8 ;
      RECT 8.95 1.7 10.3 1.95 ;
      RECT 9.9 1.65 10.3 1.95 ;
      RECT 9.9 1.05 10.15 1.95 ;
      RECT 8.1 4.9 8.6 5.2 ;
      RECT 8.2 2.3 8.5 5.2 ;
      RECT 8.1 2.3 8.6 2.6 ;
      RECT 7.1 5.05 7.35 7.25 ;
      RECT 5.45 5.05 7.35 5.3 ;
      RECT 5.45 2.35 5.7 5.3 ;
      RECT 4.4 3.6 5.7 3.9 ;
      RECT 5.45 2.35 6.45 2.6 ;
      RECT 6.05 1.65 6.45 2.6 ;
      RECT 6.05 1.65 7.35 1.9 ;
      RECT 7.1 1.05 7.35 1.9 ;
      RECT 4.7 5.8 4.95 7.25 ;
      RECT 3 5.8 3.25 7.25 ;
      RECT 3 5.8 4.95 6.05 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 4.5 2.25 4.75 2.65 ;
      RECT 3.15 2.3 4.9 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 14.95 2.25 15.45 2.55 ;
      RECT 12.95 2.25 13.45 2.55 ;
      RECT 10.1 2.95 10.6 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsr_1
