magic
tech gf180mcuC
timestamp 1660765831
<< error_p >>
rect 8 97 18 159
<< nwell >>
rect 0 97 8 159
<< metal1 >>
rect 0 147 8 159
rect 0 36 8 48
<< labels >>
rlabel metal1 4 153 4 153 3 VDD
rlabel metal1 7 41 7 41 1 GND
<< end >>
