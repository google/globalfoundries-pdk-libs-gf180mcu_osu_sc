# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffn_1 0 0 ;
  SIZE 14.25 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 14.25 8.1 ;
        RECT 12.55 5.45 12.8 8.1 ;
        RECT 9.95 5.45 10.35 8.1 ;
        RECT 7.25 6.2 7.5 8.1 ;
        RECT 4.45 5.45 4.7 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.25 0.6 ;
        RECT 12.55 0 12.8 1.8 ;
        RECT 9.95 0 10.35 1.45 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 4.45 0 4.7 1.4 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9.5 2.85 10 3.15 ;
        RECT 9.6 2.75 9.9 3.25 ;
      LAYER MET2 ;
        RECT 9.5 2.85 10 3.15 ;
        RECT 9.55 2.8 9.95 3.2 ;
      LAYER VIA12 ;
        RECT 9.62 2.87 9.88 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.5 2.4 3.8 ;
      LAYER MET2 ;
        RECT 1.75 3.5 2.55 3.8 ;
        RECT 1.9 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.02 3.52 2.28 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.4 4.8 13.9 5.15 ;
        RECT 13.4 4.75 13.85 5.15 ;
        RECT 13.4 0.95 13.65 7.15 ;
      LAYER MET2 ;
        RECT 13.4 4.8 13.9 5.1 ;
        RECT 13.45 4.75 13.85 5.15 ;
      LAYER VIA12 ;
        RECT 13.52 4.82 13.78 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.7 4.15 13.15 4.45 ;
        RECT 12.8 2.05 13.05 4.45 ;
        RECT 11.7 2.05 13.05 2.3 ;
        RECT 11.7 4.15 11.95 7.15 ;
        RECT 11.7 0.95 11.95 2.3 ;
      LAYER MET2 ;
        RECT 12.65 4.15 13.15 4.45 ;
        RECT 12.7 4.1 13.1 4.5 ;
      LAYER VIA12 ;
        RECT 12.77 4.17 13.03 4.43 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 6.75 4.75 7.15 5.15 ;
      RECT 6.7 4.8 11.15 5.1 ;
      RECT 10.85 2.85 11.15 5.1 ;
      RECT 11.95 2.8 12.35 3.2 ;
      RECT 10.85 2.85 12.4 3.15 ;
      RECT 10.25 1.65 10.65 2.05 ;
      RECT 9.5 1.7 10.7 2 ;
      RECT 5.8 1.5 6.2 1.9 ;
      RECT 5.75 1.55 9.9 1.85 ;
      RECT 5.75 1.65 10.65 1.85 ;
      RECT 8.9 4.1 9.3 4.5 ;
      RECT 7.7 4.1 8.1 4.5 ;
      RECT 6.05 4.1 6.55 4.5 ;
      RECT 3.25 4.1 3.7 4.5 ;
      RECT 3.25 4.15 9.35 4.45 ;
      RECT 8.05 2.8 8.45 3.2 ;
      RECT 6.1 2.8 6.5 3.2 ;
      RECT 6.05 2.85 8.55 3.15 ;
      RECT 6.8 3.45 7.2 3.85 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.1 2.15 4.5 2.55 ;
      RECT 0.45 2.15 0.85 2.55 ;
      RECT 0.4 2.2 4.55 2.5 ;
    LAYER VIA12 ;
      RECT 12.02 2.87 12.28 3.13 ;
      RECT 10.32 1.72 10.58 1.98 ;
      RECT 8.97 4.17 9.23 4.43 ;
      RECT 8.12 2.87 8.38 3.13 ;
      RECT 7.77 4.17 8.03 4.43 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.82 4.82 7.08 5.08 ;
      RECT 6.17 2.87 6.43 3.13 ;
      RECT 6.17 4.17 6.43 4.43 ;
      RECT 5.87 1.57 6.13 1.83 ;
      RECT 4.17 2.22 4.43 2.48 ;
      RECT 3.37 4.17 3.63 4.43 ;
      RECT 0.52 2.22 0.78 2.48 ;
    LAYER MET1 ;
      RECT 10.95 0.95 11.2 7.15 ;
      RECT 10.95 2.85 12.4 3.15 ;
      RECT 10.3 1.7 10.6 5.2 ;
      RECT 10.2 4.8 10.7 5.1 ;
      RECT 10.2 1.7 10.7 2 ;
      RECT 9.1 5.45 9.35 7.15 ;
      RECT 8.95 1.6 9.25 5.7 ;
      RECT 9.1 0.95 9.35 1.85 ;
      RECT 8.1 4.75 8.35 7.15 ;
      RECT 8.1 4.75 8.7 5 ;
      RECT 8.4 3.55 8.7 5 ;
      RECT 8.1 2.75 8.4 3.8 ;
      RECT 8.1 0.95 8.35 3.8 ;
      RECT 6.7 4.8 7.2 5.1 ;
      RECT 6.8 3.5 7.1 5.1 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 5.5 4.15 6.55 4.45 ;
      RECT 5.5 2.15 5.8 4.45 ;
      RECT 5.4 2.15 5.9 2.45 ;
      RECT 5.85 5.95 6.1 7.15 ;
      RECT 4.95 5.95 6.1 6.2 ;
      RECT 4.95 3.45 5.2 6.2 ;
      RECT 4.9 1.6 5.15 3.7 ;
      RECT 4.9 1.6 6.25 1.85 ;
      RECT 5.85 1.55 6.25 1.85 ;
      RECT 5.85 0.95 6.1 1.85 ;
      RECT 4.05 4.8 4.55 5.1 ;
      RECT 4.15 2.2 4.45 5.1 ;
      RECT 4.05 2.2 4.55 2.5 ;
      RECT 2.6 4.15 3.75 4.45 ;
      RECT 3.35 2.2 3.65 4.45 ;
      RECT 3.25 2.2 3.75 2.5 ;
      RECT 3.05 4.95 3.3 7.15 ;
      RECT 1.4 4.95 3.3 5.2 ;
      RECT 1.4 2.25 1.65 5.2 ;
      RECT 1.05 4.15 1.65 4.45 ;
      RECT 1.4 2.25 2.4 2.5 ;
      RECT 2 1.55 2.4 2.5 ;
      RECT 2 1.55 3.3 1.8 ;
      RECT 3.05 0.95 3.3 1.8 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.5 2.1 0.8 2.6 ;
      RECT 7.65 4.15 8.15 4.45 ;
      RECT 6.05 2.85 6.55 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffn_1
