* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__addf_1 A B CI S CO VDD VSS
X0 a_9_70# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_110_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 S a_161_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 S a_161_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 a_195_19# B a_178_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_178_19# A a_161_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_195_70# B a_178_70# VDD pmos_3p3 w=1.7u l=0.3u
X7 a_110_19# CI VSS VSS nmos_3p3 w=0.85u l=0.3u
X8 a_178_70# A a_161_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_59_19# CI a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS B a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_110_70# CI VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS A a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_59_19# CI a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X14 VDD B a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X15 CO a_59_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X16 VDD A a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS CI a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 CO a_59_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X19 VDD CI a_195_70# VDD pmos_3p3 w=1.7u l=0.3u
X20 VSS A a_76_19# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_161_19# a_59_19# a_110_19# VSS nmos_3p3 w=0.85u l=0.3u
X22 a_76_19# B a_59_19# VSS nmos_3p3 w=0.85u l=0.3u
X23 VDD A a_76_70# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_161_19# a_59_19# a_110_70# VDD pmos_3p3 w=1.7u l=0.3u
X25 a_9_19# B VSS VSS nmos_3p3 w=0.85u l=0.3u
X26 a_110_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X27 a_76_70# B a_59_19# VDD pmos_3p3 w=1.7u l=0.3u
.ends
