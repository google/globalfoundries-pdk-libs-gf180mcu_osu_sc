# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__buf_4
  CLASS CORE ;
  ORIGIN 0 0.05 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__buf_4 0 -0.05 ;
  SIZE 5.7 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.6 5.7 6.3 ;
        RECT 4.85 3.55 5.1 6.3 ;
        RECT 3.15 3.55 3.4 6.3 ;
        RECT 1.45 3.55 1.7 6.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.05 5.7 0.65 ;
        RECT 4.85 -0.05 5.1 1.85 ;
        RECT 3.15 -0.05 3.4 1.85 ;
        RECT 1.45 -0.05 1.7 1.85 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.1 2.25 1.6 2.55 ;
      LAYER Metal2 ;
        RECT 1.1 2.25 1.6 2.55 ;
        RECT 1.15 2.2 1.55 2.6 ;
      LAYER Via1 ;
        RECT 1.22 2.27 1.48 2.53 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.9 3.55 4.4 3.85 ;
        RECT 4 1 4.25 5.25 ;
        RECT 2.3 3 4.25 3.3 ;
        RECT 2.3 2.1 4.25 2.4 ;
        RECT 2.3 1 2.55 5.25 ;
      LAYER Metal2 ;
        RECT 3.9 3.5 4.4 3.9 ;
      LAYER Via1 ;
        RECT 4.02 3.57 4.28 3.83 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.6 1 0.85 5.25 ;
      RECT 0.6 3 2.05 3.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__buf_4
