* NGSPICE file created from gf180mcu_osu_sc_12T_buf_2.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 VDD a_n8_16# Y VDD pmos_3p3 w=1.7u l=0.3u
X1 Y a_n8_16# VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_n8_16# GND GND nmos_3p3 w=0.85u l=0.3u
X3 VDD A a_n8_16# VDD pmos_3p3 w=1.7u l=0.3u
X4 GND a_n8_16# Y GND nmos_3p3 w=0.85u l=0.3u
X5 GND A a_n8_16# GND nmos_3p3 w=0.85u l=0.3u
