* NGSPICE file created from gf180mcu_osu_sc_9T_mux2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y a_25_19# A GND nmos_3p3 w=0.85u l=0.3u
X1 a_25_19# Sel GND GND nmos_3p3 w=0.85u l=0.3u
X2 Y Sel A VDD pmos_3p3 w=1.7u l=0.3u
X3 a_25_19# Sel VDD VDD pmos_3p3 w=1.7u l=0.3u
X4 B Sel Y GND nmos_3p3 w=0.85u l=0.3u
X5 B a_25_19# Y VDD pmos_3p3 w=1.7u l=0.3u
