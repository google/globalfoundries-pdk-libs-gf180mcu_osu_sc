* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__dffn_1 D Q QN CLK VDD VSS
X0 a_42_70# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_125_19# a_53_38# a_114_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X3 a_161_42# a_125_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X4 a_86_70# a_53_38# a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X5 VDD a_161_42# a_148_70# VDD pmos_3p3 w=1.7u l=0.3u
X6 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 VSS a_9_19# a_86_19# VSS nmos_3p3 w=0.85u l=0.3u
X8 a_19_14# a_53_38# a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X9 a_161_42# a_125_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 VDD a_9_19# a_86_70# VDD pmos_3p3 w=1.7u l=0.3u
X11 a_19_14# a_50_59# a_42_70# VDD pmos_3p3 w=1.7u l=0.3u
X12 VSS a_19_14# a_9_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_53_38# a_50_59# VSS VSS nmos_3p3 w=0.85u l=0.3u
X14 VDD a_19_14# a_9_19# VDD pmos_3p3 w=1.7u l=0.3u
X15 VSS a_161_42# QN VSS nmos_3p3 w=0.85u l=0.3u
X16 a_53_38# a_50_59# VDD VDD pmos_3p3 w=1.7u l=0.3u
X17 VSS CLK a_50_59# VSS nmos_3p3 w=0.85u l=0.3u
X18 VDD a_161_42# QN VDD pmos_3p3 w=1.7u l=0.3u
X19 a_148_19# a_53_38# a_125_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_114_19# a_9_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X21 VDD CLK a_50_59# VDD pmos_3p3 w=1.7u l=0.3u
X22 a_148_70# a_50_59# a_125_19# VDD pmos_3p3 w=1.7u l=0.3u
X23 a_114_70# a_9_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 a_42_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X25 a_125_19# a_50_59# a_114_19# VSS nmos_3p3 w=0.85u l=0.3u
X26 a_86_19# a_50_59# a_19_14# VSS nmos_3p3 w=0.85u l=0.3u
X27 VSS a_161_42# a_148_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
