* NGSPICE file created from gf180mcu_osu_sc_9T_addh_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_19_14# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_91_19# B a_91_70# VDD pmos_3p3 w=1.7u l=0.3u
X2 GND a_19_14# a_75_19# GND nmos_3p3 w=0.85u l=0.3u
X3 VDD a_19_14# a_91_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 a_19_14# B a_42_19# GND nmos_3p3 w=0.85u l=0.3u
X5 GND a_19_14# CO GND nmos_3p3 w=0.85u l=0.3u
X6 VDD B a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X7 VDD a_19_14# CO VDD pmos_3p3 w=1.7u l=0.3u
X8 S a_91_19# GND GND nmos_3p3 w=0.85u l=0.3u
X9 a_91_19# A a_75_19# GND nmos_3p3 w=0.85u l=0.3u
X10 S a_91_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X11 a_42_19# A GND GND nmos_3p3 w=0.85u l=0.3u
X12 a_91_70# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 a_75_19# B a_91_19# GND nmos_3p3 w=0.85u l=0.3u
