# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__addh_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addh_1 0 0 ;
  SIZE 8.6 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 8.6 6.15 ;
        RECT 6.65 4.5 6.9 6.15 ;
        RECT 3.85 3.5 4.1 6.15 ;
        RECT 3.1 3.5 3.35 6.15 ;
        RECT 1.4 3.5 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 8.6 0.6 ;
        RECT 6.65 0 6.9 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 2.2 4.4 2.5 ;
        RECT 1.5 2.2 2 2.5 ;
      LAYER MET2 ;
        RECT 3.9 2.15 4.4 2.55 ;
        RECT 1.5 2.2 4.4 2.5 ;
        RECT 1.5 2.15 2 2.55 ;
      LAYER VIA12 ;
        RECT 1.62 2.22 1.88 2.48 ;
        RECT 4.02 2.22 4.28 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.2 1.9 5.5 2.4 ;
        RECT 2.35 2.15 2.85 2.45 ;
        RECT 2.35 1.55 2.85 1.85 ;
        RECT 2.45 1.55 2.75 2.45 ;
      LAYER MET2 ;
        RECT 5.15 1.95 5.55 2.35 ;
        RECT 5.2 1.55 5.5 2.4 ;
        RECT 5.15 1.55 5.5 2.35 ;
        RECT 2.35 1.55 5.5 1.85 ;
        RECT 2.4 1.5 2.8 1.9 ;
      LAYER VIA12 ;
        RECT 2.47 1.57 2.73 1.83 ;
        RECT 5.22 2.02 5.48 2.28 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 3.5 0.9 3.8 ;
        RECT 0.55 0.95 0.8 5.2 ;
      LAYER MET2 ;
        RECT 0.4 3.45 0.9 3.85 ;
      LAYER VIA12 ;
        RECT 0.52 3.52 0.78 3.78 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 7.7 2.85 8.2 3.15 ;
        RECT 7.75 2.8 8.1 3.2 ;
        RECT 7.5 3.5 8 5.2 ;
        RECT 7.75 0.95 8 5.2 ;
      LAYER MET2 ;
        RECT 7.7 2.8 8.2 3.2 ;
      LAYER VIA12 ;
        RECT 7.82 2.87 8.08 3.13 ;
    END
  END S
  OBS
    LAYER MET2 ;
      RECT 6.3 2.95 6.8 3.35 ;
      RECT 3 2.9 3.5 3.3 ;
      RECT 3 2.95 6.8 3.25 ;
    LAYER VIA12 ;
      RECT 6.42 3.02 6.68 3.28 ;
      RECT 3.12 2.97 3.38 3.23 ;
    LAYER MET1 ;
      RECT 5.55 3.5 6.05 5.2 ;
      RECT 5.55 2.75 5.8 5.2 ;
      RECT 4.7 2.75 6.05 3 ;
      RECT 5.75 2.5 6.75 2.75 ;
      RECT 4.7 1.35 4.95 3 ;
      RECT 6.5 2.2 7.25 2.5 ;
      RECT 5.55 0.85 5.8 1.45 ;
      RECT 3.85 0.85 4.1 1.45 ;
      RECT 3.85 0.85 5.8 1.1 ;
      RECT 2.25 2.95 2.5 5.2 ;
      RECT 1.05 2.95 3.5 3.25 ;
      RECT 3.1 0.95 3.35 3.25 ;
      RECT 6.3 3 6.8 3.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addh_1
