* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp9t3v3__lshifup A Y
X0 a_26_19 A VDDH VDDH pmos_3p3 w=34 l=6
X1 Y a_46_19 VDDH VDDH pmos_3p3 w=34 l=6
X2 VSS A a_46_19 VSS nmos_3p3 w=17 l=6
X3 VDDH a_56_55 a_46_19 VDDH pmos_3p3 w=34 l=6
X4 a_56_55 a_26_19 VSS VSS nmos_3p3 w=17 l=6
X5 a_56_55 a_46_19 VDDH VDDH pmos_3p3 w=34 l=6
X6 a_26_19 A VSS VSS nmos_3p3 w=17 l=6
X7 Y a_46_19 VSS VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
