# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dff_1 0 0 ;
  SIZE 13 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 13 8.1 ;
        RECT 11.3 5.45 11.55 8.1 ;
        RECT 8.85 5.45 9.1 8.1 ;
        RECT 7.25 6.2 7.5 8.1 ;
        RECT 4.45 5.45 4.7 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 13 0.6 ;
        RECT 11.3 0 11.55 1.8 ;
        RECT 8.85 0 9.1 1.45 ;
        RECT 7.25 0 7.5 1.8 ;
        RECT 4.45 0 4.7 1.4 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.65 4.15 8.15 4.45 ;
        RECT 5.5 4.15 6.55 4.45 ;
        RECT 5.4 2.15 5.9 2.45 ;
        RECT 5.5 2.15 5.8 4.45 ;
        RECT 2.6 4.15 3.75 4.45 ;
        RECT 3.25 2.2 3.75 2.5 ;
        RECT 3.35 2.2 3.65 4.45 ;
      LAYER MET2 ;
        RECT 3.25 4.15 8.15 4.45 ;
        RECT 7.7 4.1 8.1 4.5 ;
        RECT 6.05 4.1 6.55 4.5 ;
        RECT 3.25 4.1 3.7 4.5 ;
      LAYER VIA12 ;
        RECT 3.37 4.17 3.63 4.43 ;
        RECT 6.17 4.17 6.43 4.43 ;
        RECT 7.77 4.17 8.03 4.43 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.5 2.4 3.8 ;
      LAYER MET2 ;
        RECT 1.75 3.5 2.55 3.8 ;
        RECT 1.9 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.02 3.52 2.28 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.15 4.8 12.65 5.15 ;
        RECT 12.15 4.75 12.6 5.15 ;
        RECT 12.15 0.95 12.4 7.15 ;
      LAYER MET2 ;
        RECT 12.15 4.8 12.65 5.1 ;
        RECT 12.2 4.75 12.6 5.15 ;
      LAYER VIA12 ;
        RECT 12.27 4.82 12.53 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.45 4.15 11.9 4.45 ;
        RECT 11.55 2.05 11.8 4.45 ;
        RECT 10.45 2.05 11.8 2.3 ;
        RECT 10.45 4.15 10.7 7.15 ;
        RECT 10.45 0.95 10.7 2.3 ;
      LAYER MET2 ;
        RECT 11.4 4.15 11.9 4.45 ;
        RECT 11.45 4.1 11.85 4.5 ;
      LAYER VIA12 ;
        RECT 11.52 4.17 11.78 4.43 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 6.75 4.75 7.15 5.15 ;
      RECT 6.7 4.8 9.9 5.1 ;
      RECT 9.6 2.85 9.9 5.1 ;
      RECT 10.7 2.8 11.1 3.2 ;
      RECT 9.6 2.85 11.15 3.15 ;
      RECT 9 1.65 9.4 2.05 ;
      RECT 8.5 1.7 9.45 2 ;
      RECT 5.8 1.5 6.2 1.9 ;
      RECT 5.75 1.55 8.8 1.85 ;
      RECT 5.75 1.65 9.4 1.85 ;
      RECT 8.05 2.8 8.45 3.2 ;
      RECT 6.1 2.8 6.5 3.2 ;
      RECT 6.05 2.85 8.55 3.15 ;
      RECT 6.8 3.45 7.2 3.85 ;
      RECT 6.75 3.5 7.25 3.8 ;
      RECT 4.1 2.15 4.5 2.55 ;
      RECT 0.45 2.15 0.85 2.55 ;
      RECT 0.4 2.2 4.55 2.5 ;
    LAYER VIA12 ;
      RECT 10.77 2.87 11.03 3.13 ;
      RECT 9.07 1.72 9.33 1.98 ;
      RECT 8.12 2.87 8.38 3.13 ;
      RECT 6.87 3.52 7.13 3.78 ;
      RECT 6.82 4.82 7.08 5.08 ;
      RECT 6.17 2.87 6.43 3.13 ;
      RECT 5.87 1.57 6.13 1.83 ;
      RECT 4.17 2.22 4.43 2.48 ;
      RECT 0.52 2.22 0.78 2.48 ;
    LAYER MET1 ;
      RECT 9.7 0.95 9.95 7.15 ;
      RECT 9.7 2.85 11.15 3.15 ;
      RECT 9.05 1.7 9.35 3.25 ;
      RECT 8.95 2.85 9.45 3.15 ;
      RECT 8.95 1.7 9.45 2 ;
      RECT 8.1 4.75 8.35 7.15 ;
      RECT 8.1 4.75 8.9 5 ;
      RECT 8.6 3.55 8.9 5 ;
      RECT 8.1 3.55 8.9 3.8 ;
      RECT 8.1 2.75 8.4 3.8 ;
      RECT 8.1 0.95 8.35 3.8 ;
      RECT 6.7 4.8 7.2 5.1 ;
      RECT 6.8 3.45 7.1 5.1 ;
      RECT 6.75 3.5 7.3 3.8 ;
      RECT 6.8 3.45 7.2 3.8 ;
      RECT 5.85 5.95 6.1 7.15 ;
      RECT 4.95 5.95 6.1 6.2 ;
      RECT 4.95 3.45 5.2 6.2 ;
      RECT 4.9 1.6 5.15 3.7 ;
      RECT 4.9 1.6 6.25 1.85 ;
      RECT 5.85 1.55 6.25 1.85 ;
      RECT 5.85 0.95 6.1 1.85 ;
      RECT 4.05 4.8 4.55 5.1 ;
      RECT 4.15 2.2 4.45 5.1 ;
      RECT 4.05 2.2 4.55 2.5 ;
      RECT 3.05 4.95 3.3 7.15 ;
      RECT 1.4 4.95 3.3 5.2 ;
      RECT 1.4 2.25 1.65 5.2 ;
      RECT 1.05 4.15 1.65 4.45 ;
      RECT 1.4 2.25 2.4 2.5 ;
      RECT 2 1.55 2.4 2.5 ;
      RECT 2 1.55 3.3 1.8 ;
      RECT 3.05 0.95 3.3 1.8 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.5 2.1 0.8 2.6 ;
      RECT 6.05 2.85 6.55 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dff_1
