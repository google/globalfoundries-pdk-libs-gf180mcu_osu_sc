# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__addf_1 0 0 ;
  SIZE 14 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 14 6.35 ;
        RECT 12.35 4.8 12.6 6.35 ;
        RECT 10.75 4.8 11 6.35 ;
        RECT 6.5 4.8 6.75 6.35 ;
        RECT 4.8 4.8 5.05 6.35 ;
        RECT 1.4 4.8 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14 0.7 ;
        RECT 12.35 0 12.6 1.5 ;
        RECT 10.75 0 11 1.5 ;
        RECT 6.5 0 6.75 1.5 ;
        RECT 4.8 0 5.05 1.5 ;
        RECT 1.4 0 1.65 1.5 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.7 2.45 9.2 2.75 ;
        RECT 6.4 3.15 9.1 3.45 ;
        RECT 8.8 2.45 9.1 3.45 ;
        RECT 6.4 2.45 6.7 3.45 ;
        RECT 3.2 2.45 6.7 2.75 ;
        RECT 2.15 3.2 3.45 3.5 ;
        RECT 3.2 2.45 3.45 3.5 ;
        RECT 2.15 2.3 2.4 3.5 ;
        RECT 0.6 2.3 2.4 2.6 ;
      LAYER Metal2 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.85 3.7 9.95 4 ;
        RECT 9.65 3 9.95 4 ;
        RECT 5.85 3 6.15 4 ;
        RECT 3.7 3.1 6.15 3.4 ;
        RECT 1.6 3.75 4 4.05 ;
        RECT 3.7 3 4 4.05 ;
        RECT 1.6 2.85 1.9 4.05 ;
      LAYER Metal2 ;
        RECT 1.5 2.95 2 3.25 ;
        RECT 1.55 2.9 1.95 3.3 ;
      LAYER Via1 ;
        RECT 1.62 2.97 1.88 3.23 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.75 2.35 10.6 2.65 ;
        RECT 9.75 1.9 10.05 2.65 ;
        RECT 2.65 1.9 10.05 2.2 ;
        RECT 7.05 1.9 7.35 2.85 ;
        RECT 2.65 1.9 2.95 2.7 ;
      LAYER Metal2 ;
        RECT 2.55 2.3 3.05 2.6 ;
        RECT 2.6 2.25 3 2.65 ;
      LAYER Via1 ;
        RECT 2.67 2.32 2.93 2.58 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.2 3.1 13.75 3.4 ;
        RECT 13.2 3.05 13.65 3.45 ;
        RECT 13.2 1.05 13.45 5.3 ;
      LAYER Metal2 ;
        RECT 13.25 3.1 13.75 3.4 ;
        RECT 13.3 3.05 13.7 3.45 ;
      LAYER Via1 ;
        RECT 13.37 3.12 13.63 3.38 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.6 3.1 12.05 3.4 ;
        RECT 11.6 3.05 11.9 3.45 ;
        RECT 11.6 1.05 11.85 5.3 ;
      LAYER Metal2 ;
        RECT 11.55 3.1 12.05 3.4 ;
        RECT 11.6 3.05 12 3.45 ;
      LAYER Via1 ;
        RECT 11.67 3.12 11.93 3.38 ;
    END
  END S
  OBS
    LAYER Metal2 ;
      RECT 3.1 4.85 3.4 5.3 ;
      RECT 3.05 4.85 3.45 5.25 ;
      RECT 3 4.9 12.85 5.2 ;
      RECT 12.55 2.35 12.85 5.2 ;
      RECT 3.75 1.15 4.05 5.2 ;
      RECT 12.5 2.4 12.9 2.8 ;
      RECT 7.85 2.4 8.25 2.8 ;
      RECT 12.45 2.45 12.95 2.75 ;
      RECT 3.75 2.45 8.3 2.75 ;
      RECT 3.1 1.05 3.4 1.55 ;
      RECT 3.05 1.1 3.45 1.5 ;
      RECT 3.05 1.15 4.05 1.45 ;
      RECT 8.15 4.2 8.55 4.6 ;
      RECT 8.1 4.25 11.25 4.55 ;
      RECT 10.95 2.35 11.25 4.55 ;
      RECT 8.85 1.15 9.15 4.55 ;
      RECT 10.9 2.4 11.3 2.8 ;
      RECT 8.15 1.1 8.55 1.5 ;
      RECT 8.1 1.15 9.15 1.45 ;
      RECT 7.3 1.05 7.6 1.55 ;
      RECT 5.65 1.05 5.95 1.55 ;
      RECT 7.25 1.1 7.65 1.5 ;
      RECT 5.6 1.1 6 1.5 ;
      RECT 5.6 1.15 7.65 1.45 ;
      RECT 2.2 1.05 2.5 1.55 ;
      RECT 0.5 1.05 0.8 1.55 ;
      RECT 2.15 1.1 2.55 1.5 ;
      RECT 0.45 1.1 0.85 1.5 ;
      RECT 0.45 1.15 2.55 1.45 ;
    LAYER Via1 ;
      RECT 12.57 2.47 12.83 2.73 ;
      RECT 10.97 2.47 11.23 2.73 ;
      RECT 8.22 1.17 8.48 1.43 ;
      RECT 8.22 4.27 8.48 4.53 ;
      RECT 7.92 2.47 8.18 2.73 ;
      RECT 7.32 1.17 7.58 1.43 ;
      RECT 5.67 1.17 5.93 1.43 ;
      RECT 3.12 1.17 3.38 1.43 ;
      RECT 3.12 4.92 3.38 5.18 ;
      RECT 2.22 1.17 2.48 1.43 ;
      RECT 0.52 1.17 0.78 1.43 ;
    LAYER Metal1 ;
      RECT 7.35 4.3 7.6 5.3 ;
      RECT 5.65 4.3 5.9 5.3 ;
      RECT 5.65 4.3 7.6 4.55 ;
      RECT 2.25 4.3 2.5 5.3 ;
      RECT 0.55 4.3 0.8 5.3 ;
      RECT 0.55 4.3 2.5 4.55 ;
      RECT 12.45 2.45 12.95 2.75 ;
      RECT 10.85 2.45 11.35 2.75 ;
      RECT 8.1 4.25 8.6 4.55 ;
      RECT 8.2 1.05 8.5 1.55 ;
      RECT 7.8 2.45 8.3 2.75 ;
      RECT 7.3 1.05 7.6 1.55 ;
      RECT 5.65 1.05 5.95 1.55 ;
      RECT 3.1 1.05 3.4 1.55 ;
      RECT 3.1 4.8 3.4 5.3 ;
      RECT 2.2 1.05 2.5 1.55 ;
      RECT 0.5 1.05 0.8 1.55 ;
  END
END gf180mcu_osu_sc_gp9t3v3__addf_1
