* include file for sky130 models

.lib 'sky130.lib.spice' TT
