# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_1 0 0 ;
  SIZE 3.85 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.85 6.15 ;
        RECT 1.4 3.5 1.75 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.85 0.6 ;
        RECT 1.4 0 1.75 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.2 2.1 2.5 ;
      LAYER MET2 ;
        RECT 1.6 2.2 2.1 2.5 ;
        RECT 1.65 2.15 2.05 2.55 ;
      LAYER VIA12 ;
        RECT 1.72 2.22 1.98 2.48 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 1.9 2.8 2.4 ;
        RECT 0.8 2.2 1.3 2.5 ;
      LAYER MET2 ;
        RECT 2.4 1.95 2.9 2.35 ;
        RECT 2.4 1.55 2.8 2.35 ;
        RECT 0.9 1.55 2.8 1.85 ;
        RECT 0.8 2.2 1.3 2.5 ;
        RECT 0.85 2.15 1.25 2.55 ;
        RECT 0.9 1.55 1.2 2.55 ;
      LAYER VIA12 ;
        RECT 0.92 2.22 1.18 2.48 ;
        RECT 2.52 2.02 2.78 2.28 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.15 1.25 3.4 4.05 ;
        RECT 2.9 3.75 3.2 4.55 ;
        RECT 2.9 3.75 3.15 5.2 ;
        RECT 2.9 0.95 3.15 1.5 ;
      LAYER MET2 ;
        RECT 2.8 4.1 3.3 4.5 ;
      LAYER VIA12 ;
        RECT 2.92 4.17 3.18 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 0.4 3.45 0.9 3.85 ;
      RECT 0.4 3.5 2 3.8 ;
      RECT 1.7 3 2 3.8 ;
      RECT 2.4 2.95 2.9 3.35 ;
      RECT 1.7 3 2.9 3.3 ;
    LAYER VIA12 ;
      RECT 2.52 3.02 2.78 3.28 ;
      RECT 0.52 3.52 0.78 3.78 ;
    LAYER MET1 ;
      RECT 0.55 2.95 0.8 5.2 ;
      RECT 0.4 3.5 0.9 3.8 ;
      RECT 0.3 1.55 0.55 3.2 ;
      RECT 0.55 0.95 0.8 1.8 ;
      RECT 2.5 2.9 2.8 3.4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_1
