# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffrn_1 0 0 ;
  SIZE 19.25 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 19.25 8.3 ;
        RECT 17.6 5.55 17.85 8.3 ;
        RECT 14.6 5.55 14.85 8.3 ;
        RECT 13.4 5.55 13.65 8.3 ;
        RECT 10.75 6.3 11 8.3 ;
        RECT 7.95 5.55 8.2 8.3 ;
        RECT 4.9 5.55 5.15 8.3 ;
        RECT 3.55 5.55 3.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 19.25 0.7 ;
        RECT 17.6 0 17.85 1.9 ;
        RECT 15.85 0 16.1 1.9 ;
        RECT 14.15 0 14.4 1.9 ;
        RECT 13.4 0 13.65 1.9 ;
        RECT 10.75 0 11 1.9 ;
        RECT 7.95 0 8.2 1.5 ;
        RECT 4.9 0 5.15 1.9 ;
        RECT 4 0 4.25 1.9 ;
        RECT 2.3 0 2.55 1.9 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 13.15 2.95 13.65 3.25 ;
      LAYER Metal2 ;
        RECT 13.15 2.9 13.65 3.3 ;
      LAYER Via1 ;
        RECT 13.27 2.97 13.53 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.4 3.6 5.9 3.9 ;
      LAYER Metal2 ;
        RECT 5.4 3.55 5.9 3.95 ;
      LAYER Via1 ;
        RECT 5.52 3.62 5.78 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 18.45 4.9 18.95 5.25 ;
        RECT 18.45 4.85 18.9 5.25 ;
        RECT 18.45 1.05 18.7 7.25 ;
      LAYER Metal2 ;
        RECT 18.45 4.9 18.95 5.2 ;
        RECT 18.5 4.85 18.9 5.25 ;
      LAYER Via1 ;
        RECT 18.57 4.92 18.83 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 16.75 4.25 18.2 4.55 ;
        RECT 17.85 2.15 18.1 4.55 ;
        RECT 16.75 2.15 18.1 2.4 ;
        RECT 16.75 4.25 17 7.25 ;
        RECT 16.75 1.05 17 2.4 ;
      LAYER Metal2 ;
        RECT 17.7 4.25 18.2 4.55 ;
        RECT 17.75 4.2 18.15 4.6 ;
      LAYER Via1 ;
        RECT 17.82 4.27 18.08 4.53 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 4.9 1.05 5.2 ;
      LAYER Metal2 ;
        RECT 0.55 4.85 1.05 5.25 ;
      LAYER Via1 ;
        RECT 0.67 4.92 0.93 5.18 ;
    END
  END RN
  OBS
    LAYER Metal2 ;
      RECT 17 2.9 17.4 3.3 ;
      RECT 16.65 2.95 17.45 3.25 ;
      RECT 2.65 3.55 3.15 3.95 ;
      RECT 2.75 1 3.05 3.95 ;
      RECT 1.3 2.25 1.8 2.65 ;
      RECT 15.4 2.2 16 2.6 ;
      RECT 1.3 2.3 3.05 2.6 ;
      RECT 15.4 1 15.7 2.6 ;
      RECT 2.75 1 15.7 1.3 ;
      RECT 14.05 2.2 14.55 2.6 ;
      RECT 14.05 1.65 14.45 2.6 ;
      RECT 9.3 1.6 9.7 2 ;
      RECT 9.25 1.65 14.45 1.95 ;
      RECT 14.1 4.85 14.5 5.25 ;
      RECT 10.25 4.85 10.65 5.25 ;
      RECT 10.2 4.9 14.55 5.2 ;
      RECT 12.45 4.2 12.9 4.6 ;
      RECT 11.2 4.2 11.6 4.6 ;
      RECT 9.55 4.2 10.05 4.6 ;
      RECT 6.75 4.2 7.2 4.6 ;
      RECT 6.75 4.25 12.9 4.55 ;
      RECT 11.55 2.9 11.95 3.3 ;
      RECT 9.6 2.9 10 3.3 ;
      RECT 9.55 2.95 12.05 3.25 ;
      RECT 10.3 3.55 10.7 3.95 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 7.6 2.25 8 2.65 ;
      RECT 3.85 2.25 4.35 2.65 ;
      RECT 3.85 2.3 8.05 2.6 ;
      RECT 15.9 4.85 16.4 5.25 ;
    LAYER Via1 ;
      RECT 17.07 2.97 17.33 3.23 ;
      RECT 16.02 4.92 16.28 5.18 ;
      RECT 15.62 2.27 15.88 2.53 ;
      RECT 14.17 2.27 14.43 2.53 ;
      RECT 14.17 4.92 14.43 5.18 ;
      RECT 12.52 4.27 12.78 4.53 ;
      RECT 11.62 2.97 11.88 3.23 ;
      RECT 11.27 4.27 11.53 4.53 ;
      RECT 10.37 3.62 10.63 3.88 ;
      RECT 10.32 4.92 10.58 5.18 ;
      RECT 9.67 2.97 9.93 3.23 ;
      RECT 9.67 4.27 9.93 4.53 ;
      RECT 9.37 1.67 9.63 1.93 ;
      RECT 7.67 2.32 7.93 2.58 ;
      RECT 6.87 4.27 7.13 4.53 ;
      RECT 3.97 2.32 4.23 2.58 ;
      RECT 2.77 3.62 3.03 3.88 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 16 2.95 16.25 7.25 ;
      RECT 14.15 4.8 14.45 5.3 ;
      RECT 14.15 4.9 16.4 5.2 ;
      RECT 15 2.95 17.45 3.25 ;
      RECT 15 1.05 15.25 3.25 ;
      RECT 12.55 1.05 12.8 7.25 ;
      RECT 12.4 4.25 12.9 4.55 ;
      RECT 11.6 4.85 11.85 7.25 ;
      RECT 11.6 4.85 12.15 5.1 ;
      RECT 11.9 3.65 12.15 5.1 ;
      RECT 11.6 2.85 11.9 3.9 ;
      RECT 11.6 1.05 11.85 3.9 ;
      RECT 10.2 4.9 10.7 5.2 ;
      RECT 10.3 3.6 10.6 5.2 ;
      RECT 10.25 3.6 10.75 3.9 ;
      RECT 9 4.25 10.05 4.55 ;
      RECT 9 2.25 9.3 4.55 ;
      RECT 8.9 2.25 9.4 2.55 ;
      RECT 9.35 6.05 9.6 7.25 ;
      RECT 8.45 6.05 9.6 6.3 ;
      RECT 8.45 3.55 8.7 6.3 ;
      RECT 8.4 1.7 8.65 3.8 ;
      RECT 8.4 1.7 9.75 1.95 ;
      RECT 9.35 1.65 9.75 1.95 ;
      RECT 9.35 1.05 9.6 1.95 ;
      RECT 7.55 4.9 8.05 5.2 ;
      RECT 7.65 2.3 7.95 5.2 ;
      RECT 7.55 2.3 8.05 2.6 ;
      RECT 6.1 4.25 7.25 4.55 ;
      RECT 6.85 2.3 7.15 4.55 ;
      RECT 6.75 2.3 7.25 2.6 ;
      RECT 6.55 5.05 6.8 7.25 ;
      RECT 4.9 5.05 6.8 5.3 ;
      RECT 4.9 2.35 5.15 5.3 ;
      RECT 3.85 4.25 5.15 4.55 ;
      RECT 4.9 2.35 5.9 2.6 ;
      RECT 5.5 1.65 5.9 2.6 ;
      RECT 5.5 1.65 6.8 1.9 ;
      RECT 6.55 1.05 6.8 1.9 ;
      RECT 2.15 2.6 2.4 7.25 ;
      RECT 2.15 2.6 3.4 2.85 ;
      RECT 3.15 1.05 3.4 2.85 ;
      RECT 3.95 2.25 4.2 2.65 ;
      RECT 3 2.3 4.35 2.6 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.3 2.3 1.8 2.6 ;
      RECT 1.4 2.25 1.7 2.6 ;
      RECT 15.5 2.25 16 2.55 ;
      RECT 14.05 2.25 14.55 2.55 ;
      RECT 11.15 4.25 11.65 4.55 ;
      RECT 9.55 2.95 10.05 3.25 ;
      RECT 2.65 3.6 3.15 3.9 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffrn_1
