# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffsn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffsn_1 0 0 ;
  SIZE 15.5 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15.5 8.1 ;
        RECT 13.8 5.45 14.05 8.1 ;
        RECT 11.35 6.7 11.6 8.1 ;
        RECT 8.9 6.2 9.15 8.1 ;
        RECT 6.1 5.45 6.35 8.1 ;
        RECT 3.05 5.45 3.3 8.1 ;
        RECT 1.45 6.2 1.7 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.5 0.6 ;
        RECT 13.8 0 14.05 1.8 ;
        RECT 10.65 0 10.9 1.8 ;
        RECT 8.9 0 9.15 1.8 ;
        RECT 6.1 0 6.35 1.4 ;
        RECT 3.05 0 3.3 1.8 ;
        RECT 2.15 0 2.4 1.8 ;
    END
  END VSS
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9.3 4.15 9.8 4.45 ;
        RECT 7.15 4.15 8.2 4.45 ;
        RECT 7.05 2.15 7.55 2.45 ;
        RECT 7.15 2.15 7.45 4.45 ;
        RECT 4.25 4.15 5.4 4.45 ;
        RECT 4.9 2.2 5.4 2.5 ;
        RECT 5 2.2 5.3 4.45 ;
      LAYER MET2 ;
        RECT 4.9 4.15 9.8 4.45 ;
        RECT 9.35 4.1 9.75 4.5 ;
        RECT 7.7 4.1 8.2 4.5 ;
        RECT 4.9 4.1 5.35 4.5 ;
      LAYER VIA12 ;
        RECT 5.02 4.17 5.28 4.43 ;
        RECT 7.82 4.17 8.08 4.43 ;
        RECT 9.42 4.17 9.68 4.43 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.55 3.5 4.05 3.8 ;
      LAYER MET2 ;
        RECT 3.55 3.45 4.05 3.85 ;
      LAYER VIA12 ;
        RECT 3.67 3.52 3.93 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 14.65 4.8 15.15 5.15 ;
        RECT 14.65 4.75 15.1 5.15 ;
        RECT 14.65 0.95 14.9 7.15 ;
      LAYER MET2 ;
        RECT 14.65 4.8 15.15 5.1 ;
        RECT 14.7 4.75 15.1 5.15 ;
      LAYER VIA12 ;
        RECT 14.77 4.82 15.03 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.95 4.15 14.4 4.45 ;
        RECT 14.05 2.05 14.3 4.45 ;
        RECT 12.95 2.05 14.3 2.3 ;
        RECT 12.95 4.15 13.2 7.15 ;
        RECT 12.95 0.95 13.2 2.3 ;
      LAYER MET2 ;
        RECT 13.9 4.15 14.4 4.45 ;
        RECT 13.95 4.1 14.35 4.5 ;
      LAYER VIA12 ;
        RECT 14.02 4.17 14.28 4.43 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.55 4.15 12.05 4.45 ;
        RECT 5.7 4.8 6.2 5.1 ;
        RECT 5.7 2.2 6.2 2.5 ;
        RECT 5.8 2.2 6.1 5.1 ;
        RECT 2.3 5.7 2.55 7.15 ;
        RECT 0.75 2.2 2.5 2.5 ;
        RECT 2.1 2.15 2.35 2.55 ;
        RECT 0.6 5.7 2.55 5.95 ;
        RECT 0.75 4.15 1.5 4.45 ;
        RECT 0.75 0.95 1 5.95 ;
        RECT 0.6 5.7 0.85 7.15 ;
      LAYER MET2 ;
        RECT 11.55 4.1 12.05 4.5 ;
        RECT 1.1 5.45 11.95 5.75 ;
        RECT 11.65 4.1 11.95 5.75 ;
        RECT 1 4.1 1.5 4.5 ;
        RECT 1.1 4.1 1.4 5.75 ;
        RECT 2 2.2 6.2 2.5 ;
        RECT 5.75 2.15 6.15 2.55 ;
        RECT 2 2.15 2.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.12 4.17 1.38 4.43 ;
        RECT 2.12 2.22 2.38 2.48 ;
        RECT 5.82 2.22 6.08 2.48 ;
        RECT 11.67 4.17 11.93 4.43 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 13.2 2.8 13.6 3.2 ;
      RECT 12.85 2.85 13.65 3.15 ;
      RECT 10.55 2.1 11.05 2.5 ;
      RECT 10.55 1.55 10.95 2.5 ;
      RECT 7.45 1.5 7.85 1.9 ;
      RECT 7.4 1.55 10.95 1.85 ;
      RECT 10.6 4.75 11 5.15 ;
      RECT 8.4 4.75 8.8 5.15 ;
      RECT 8.35 4.8 11.05 5.1 ;
      RECT 9.7 2.8 10.1 3.2 ;
      RECT 7.75 2.8 8.15 3.2 ;
      RECT 7.7 2.85 10.2 3.15 ;
      RECT 8.45 3.45 8.85 3.85 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 12.25 4.75 12.75 5.15 ;
      RECT 2 3.45 2.5 3.85 ;
    LAYER VIA12 ;
      RECT 13.27 2.87 13.53 3.13 ;
      RECT 12.37 4.82 12.63 5.08 ;
      RECT 10.67 2.17 10.93 2.43 ;
      RECT 10.67 4.82 10.93 5.08 ;
      RECT 9.77 2.87 10.03 3.13 ;
      RECT 8.52 3.52 8.78 3.78 ;
      RECT 8.47 4.82 8.73 5.08 ;
      RECT 7.82 2.87 8.08 3.13 ;
      RECT 7.52 1.57 7.78 1.83 ;
      RECT 2.12 3.52 2.38 3.78 ;
    LAYER MET1 ;
      RECT 12.35 2.85 12.65 5.2 ;
      RECT 10.65 4.7 10.95 5.2 ;
      RECT 10.65 4.8 12.65 5.1 ;
      RECT 12.05 2.85 13.65 3.15 ;
      RECT 12.05 0.95 12.3 3.15 ;
      RECT 12.2 6.2 12.45 7.15 ;
      RECT 10.5 6.2 10.75 7.15 ;
      RECT 10.5 6.2 12.45 6.45 ;
      RECT 9.75 4.75 10 7.15 ;
      RECT 9.75 4.75 10.3 5 ;
      RECT 10.05 3.55 10.3 5 ;
      RECT 9.75 2.75 10.05 3.8 ;
      RECT 9.75 0.95 10 3.8 ;
      RECT 8.35 4.8 8.85 5.1 ;
      RECT 8.45 3.5 8.75 5.1 ;
      RECT 8.4 3.5 8.9 3.8 ;
      RECT 7.5 5.95 7.75 7.15 ;
      RECT 6.6 5.95 7.75 6.2 ;
      RECT 6.6 3.45 6.85 6.2 ;
      RECT 6.55 1.6 6.8 3.7 ;
      RECT 6.55 1.6 7.9 1.85 ;
      RECT 7.5 1.55 7.9 1.85 ;
      RECT 7.5 0.95 7.75 1.85 ;
      RECT 4.7 4.95 4.95 7.15 ;
      RECT 3.05 4.95 4.95 5.2 ;
      RECT 3.05 2.25 3.3 5.2 ;
      RECT 2 3.5 3.3 3.8 ;
      RECT 3.05 2.25 4.05 2.5 ;
      RECT 3.65 1.55 4.05 2.5 ;
      RECT 3.65 1.55 4.95 1.8 ;
      RECT 4.7 0.95 4.95 1.8 ;
      RECT 10.55 2.15 11.05 2.45 ;
      RECT 7.7 2.85 8.2 3.15 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffsn_1
