# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_buf_2
  CLASS CORE ;
  ORIGIN 0.85 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_buf_2 -0.85 -0.15 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.2 4 0.7 4.3 ;
      LAYER MET2 ;
        RECT 0.2 4 0.7 4.3 ;
        RECT 0.25 3.95 0.65 4.35 ;
      LAYER VIA12 ;
        RECT 0.32 4.02 0.58 4.28 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -0.85 7.35 3.05 7.95 ;
        RECT 2.25 5.3 2.5 7.95 ;
        RECT 0.55 5.3 0.8 7.95 ;
      LAYER MET2 ;
        RECT 0.8 7.4 1.3 7.7 ;
        RECT 0.85 7.35 1.25 7.75 ;
        RECT -0.4 7.4 0.1 7.7 ;
        RECT -0.35 7.35 0.05 7.75 ;
      LAYER VIA12 ;
        RECT -0.28 7.42 -0.02 7.68 ;
        RECT 0.92 7.42 1.18 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -0.85 -0.15 3.05 0.45 ;
        RECT 2.25 -0.15 2.5 1.65 ;
        RECT 0.55 -0.15 0.8 1.65 ;
      LAYER MET2 ;
        RECT 0.8 0.1 1.3 0.4 ;
        RECT 0.85 0.05 1.25 0.45 ;
        RECT -0.4 0.1 0.1 0.4 ;
        RECT -0.35 0.05 0.05 0.45 ;
      LAYER VIA12 ;
        RECT -0.28 0.12 -0.02 0.38 ;
        RECT 0.92 0.12 1.18 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 4.7 1.8 5 ;
        RECT 1.4 0.8 1.65 7 ;
      LAYER MET2 ;
        RECT 1.3 4.65 1.8 5.05 ;
      LAYER VIA12 ;
        RECT 1.42 4.72 1.68 4.98 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT -0.3 0.8 -0.05 7 ;
      RECT -0.3 2.75 1.15 3.05 ;
  END
END gf180mcu_osu_sc_12T_buf_2
