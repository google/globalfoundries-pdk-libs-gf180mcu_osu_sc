magic
tech gf180mcuC
timestamp 1661533174
<< nwell >>
rect 0 97 128 159
<< nmos >>
rect 19 55 25 72
rect 36 55 42 72
rect 49 55 55 72
rect 72 55 78 72
rect 85 55 91 72
rect 102 55 108 72
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 49 106 55 140
rect 72 106 78 140
rect 85 106 91 140
rect 102 106 108 140
<< ndiff >>
rect 58 72 68 73
rect 9 70 19 72
rect 9 57 11 70
rect 16 57 19 70
rect 9 55 19 57
rect 25 70 36 72
rect 25 57 28 70
rect 33 57 36 70
rect 25 55 36 57
rect 42 55 49 72
rect 55 71 72 72
rect 55 57 61 71
rect 66 57 72 71
rect 55 55 72 57
rect 78 55 85 72
rect 91 70 102 72
rect 91 57 94 70
rect 99 57 102 70
rect 91 55 102 57
rect 108 70 118 72
rect 108 57 111 70
rect 116 57 118 70
rect 108 55 118 57
<< pdiff >>
rect 9 138 19 140
rect 9 130 11 138
rect 16 130 19 138
rect 9 106 19 130
rect 25 138 36 140
rect 25 130 28 138
rect 33 130 36 138
rect 25 106 36 130
rect 42 106 49 140
rect 55 138 72 140
rect 55 130 61 138
rect 66 130 72 138
rect 55 106 72 130
rect 78 106 85 140
rect 91 138 102 140
rect 91 130 94 138
rect 99 130 102 138
rect 91 106 102 130
rect 108 138 118 140
rect 108 130 111 138
rect 116 130 118 138
rect 108 106 118 130
<< ndiffc >>
rect 11 57 16 70
rect 28 57 33 70
rect 61 57 66 71
rect 94 57 99 70
rect 111 57 116 70
<< pdiffc >>
rect 11 130 16 138
rect 28 130 33 138
rect 61 130 66 138
rect 94 130 99 138
rect 111 130 116 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
rect 57 46 66 48
rect 57 41 59 46
rect 64 41 66 46
rect 57 39 66 41
rect 81 46 90 48
rect 81 41 83 46
rect 88 41 90 46
rect 81 39 90 41
rect 105 46 114 48
rect 105 41 107 46
rect 112 41 114 46
rect 105 39 114 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
rect 81 154 90 156
rect 81 149 83 154
rect 88 149 90 154
rect 81 147 90 149
rect 105 154 114 156
rect 105 149 107 154
rect 112 149 114 154
rect 105 147 114 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
rect 59 41 64 46
rect 83 41 88 46
rect 107 41 112 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
rect 83 149 88 154
rect 107 149 112 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 49 140 55 145
rect 72 140 78 145
rect 85 140 91 145
rect 102 140 108 145
rect 19 88 25 106
rect 36 104 42 106
rect 31 102 42 104
rect 31 96 33 102
rect 39 96 42 102
rect 31 94 42 96
rect 49 104 55 106
rect 72 104 78 106
rect 85 104 91 106
rect 102 104 108 106
rect 49 102 63 104
rect 49 96 55 102
rect 61 96 63 102
rect 49 94 63 96
rect 70 102 80 104
rect 70 96 72 102
rect 78 96 80 102
rect 85 99 108 104
rect 70 94 80 96
rect 19 86 35 88
rect 19 80 27 86
rect 33 85 35 86
rect 33 80 42 85
rect 19 78 42 80
rect 19 72 25 78
rect 36 72 42 78
rect 49 72 55 94
rect 102 88 108 99
rect 60 86 70 88
rect 91 86 108 88
rect 60 80 62 86
rect 68 80 78 86
rect 91 83 93 86
rect 60 78 78 80
rect 72 72 78 78
rect 85 80 93 83
rect 99 80 108 86
rect 85 78 108 80
rect 85 72 91 78
rect 102 72 108 78
rect 19 50 25 55
rect 36 50 42 55
rect 49 50 55 55
rect 72 50 78 55
rect 85 50 91 55
rect 102 50 108 55
<< polycontact >>
rect 33 96 39 102
rect 55 96 61 102
rect 72 96 78 102
rect 27 80 33 86
rect 62 80 68 86
rect 93 80 99 86
<< metal1 >>
rect 0 154 128 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 83 154
rect 89 148 107 154
rect 113 148 128 154
rect 0 147 128 148
rect 11 138 16 140
rect 11 102 16 130
rect 28 138 33 147
rect 61 138 66 140
rect 28 128 33 130
rect 60 130 61 131
rect 60 125 66 130
rect 94 138 99 147
rect 94 128 99 130
rect 111 138 116 140
rect 60 117 66 119
rect 111 112 116 130
rect 55 107 116 112
rect 55 102 61 107
rect 11 96 33 102
rect 39 96 48 102
rect 11 70 16 96
rect 42 86 48 96
rect 70 96 72 102
rect 78 96 80 102
rect 55 94 61 96
rect 25 80 27 86
rect 33 80 35 86
rect 42 80 62 86
rect 68 80 70 86
rect 91 80 93 86
rect 99 80 101 86
rect 60 73 66 75
rect 11 55 16 57
rect 28 70 33 72
rect 60 64 61 67
rect 28 48 33 57
rect 61 55 66 57
rect 94 70 99 72
rect 94 48 99 57
rect 111 70 116 107
rect 111 55 116 57
rect 0 47 128 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 59 47
rect 65 41 83 47
rect 89 41 107 47
rect 113 41 128 47
rect 0 36 128 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 83 149 88 154
rect 88 149 89 154
rect 83 148 89 149
rect 107 149 112 154
rect 112 149 113 154
rect 107 148 113 149
rect 60 119 66 125
rect 72 96 78 102
rect 27 80 33 86
rect 93 80 99 86
rect 60 71 66 73
rect 60 67 61 71
rect 61 67 66 71
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
rect 59 46 65 47
rect 59 41 64 46
rect 64 41 65 46
rect 83 46 89 47
rect 83 41 88 46
rect 88 41 89 46
rect 107 46 113 47
rect 107 41 112 46
rect 112 41 113 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 81 148 83 154
rect 89 148 91 154
rect 105 148 107 154
rect 113 148 115 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 60 126 66 131
rect 59 125 67 126
rect 59 119 60 125
rect 66 119 67 125
rect 59 118 67 119
rect 59 117 66 118
rect 27 87 33 88
rect 26 86 34 87
rect 26 80 27 86
rect 33 80 34 86
rect 26 79 34 80
rect 27 60 33 79
rect 59 74 65 117
rect 72 103 79 104
rect 71 102 80 103
rect 71 96 72 102
rect 78 96 80 102
rect 71 95 80 96
rect 72 94 80 95
rect 58 73 68 74
rect 58 67 60 73
rect 66 67 68 73
rect 58 66 68 67
rect 74 60 80 94
rect 93 87 99 88
rect 92 86 100 87
rect 91 80 93 86
rect 99 80 101 86
rect 92 79 100 80
rect 93 78 99 79
rect 27 54 80 60
rect 10 47 18 48
rect 34 47 42 48
rect 58 47 66 48
rect 82 47 90 48
rect 106 47 114 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 57 41 59 47
rect 65 41 67 47
rect 81 41 83 47
rect 89 41 91 47
rect 105 41 107 47
rect 113 41 115 47
rect 10 40 18 41
rect 34 40 42 41
rect 58 40 66 41
rect 82 40 90 41
rect 106 40 114 41
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 14 44 14 44 1 GND
rlabel metal2 30 83 30 83 1 A
port 1 n
rlabel metal2 96 83 96 83 1 B
port 4 n
rlabel metal2 63 121 63 121 1 Y
port 3 n
<< end >>
