# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_aoi22_1 0 0 ;
  SIZE 5.35 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 5.35 8.1 ;
        RECT 1.4 6.2 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 5.35 0.6 ;
        RECT 3.5 0 3.75 1.8 ;
        RECT 0.7 0 0.95 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.5 1.1 3.8 ;
      LAYER MET2 ;
        RECT 0.6 3.45 1.1 3.85 ;
      LAYER VIA12 ;
        RECT 0.72 3.52 0.98 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 4.15 2.1 4.45 ;
      LAYER MET2 ;
        RECT 1.6 4.1 2.1 4.5 ;
      LAYER VIA12 ;
        RECT 1.72 4.17 1.98 4.43 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 3.5 2.85 3.8 ;
      LAYER MET2 ;
        RECT 2.35 3.45 2.85 3.85 ;
      LAYER VIA12 ;
        RECT 2.47 3.52 2.73 3.78 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.3 4.15 3.8 4.45 ;
      LAYER MET2 ;
        RECT 3.3 4.1 3.8 4.5 ;
      LAYER VIA12 ;
        RECT 3.42 4.17 3.68 4.43 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.3 4.8 4.8 5.1 ;
        RECT 4.45 6 4.75 6.5 ;
        RECT 4.45 4.8 4.7 6.5 ;
        RECT 4.4 3 4.65 5.1 ;
        RECT 2.1 3 4.65 3.25 ;
        RECT 2.1 0.95 2.35 3.25 ;
        RECT 3 6.1 3.5 6.4 ;
        RECT 3.1 6.1 3.35 7.15 ;
      LAYER MET2 ;
        RECT 4.35 6.05 4.85 6.45 ;
        RECT 3 6.1 4.85 6.4 ;
        RECT 3 6.05 3.5 6.45 ;
        RECT 4.3 4.75 4.8 5.15 ;
      LAYER VIA12 ;
        RECT 3.12 6.12 3.38 6.38 ;
        RECT 4.42 4.82 4.68 5.08 ;
        RECT 4.47 6.12 4.73 6.38 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.95 5.6 4.2 7.15 ;
      RECT 2.25 5.6 2.5 7.15 ;
      RECT 0.55 5.6 0.8 7.15 ;
      RECT 0.55 5.6 4.2 5.85 ;
  END
END gf180mcu_osu_sc_12T_aoi22_1
