# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffsr_1 0 0 ;
  SIZE 20.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 20.5 6.15 ;
        RECT 18.8 4.05 19.05 6.15 ;
        RECT 15.5 4.25 15.75 6.15 ;
        RECT 12.9 4.75 13.15 6.15 ;
        RECT 9.3 4.1 9.55 6.15 ;
        RECT 5.7 4.75 5.95 6.15 ;
        RECT 3.85 4.25 4.1 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 20.5 0.6 ;
        RECT 18.8 0 19.05 1.6 ;
        RECT 17.05 0 17.3 1.4 ;
        RECT 14.8 0 15.05 1.8 ;
        RECT 12.9 0 13.15 1.7 ;
        RECT 9.3 0 9.55 1.4 ;
        RECT 5.7 0 5.95 1.5 ;
        RECT 4.55 0 4.8 1.45 ;
        RECT 2.3 0 2.55 1.4 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 13.3 2.85 13.8 3.15 ;
        RECT 6.8 3 13.7 3.3 ;
        RECT 10.25 2.2 10.75 2.45 ;
        RECT 10.35 2.2 10.65 3.3 ;
        RECT 8.1 2.15 8.6 2.45 ;
        RECT 8.2 2.15 8.5 3.3 ;
      LAYER MET2 ;
        RECT 13.3 2.85 13.8 3.15 ;
        RECT 13.35 2.8 13.75 3.2 ;
      LAYER VIA12 ;
        RECT 13.42 2.87 13.68 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.05 2.85 6.55 3.15 ;
      LAYER MET2 ;
        RECT 6 2.85 6.6 3.15 ;
        RECT 6.05 2.8 6.55 3.2 ;
      LAYER VIA12 ;
        RECT 6.17 2.87 6.43 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 19.65 0.95 19.9 5.2 ;
        RECT 19.6 4.05 19.9 4.55 ;
      LAYER MET2 ;
        RECT 19.5 4.15 20 4.45 ;
        RECT 19.55 4.1 19.95 4.5 ;
      LAYER VIA12 ;
        RECT 19.62 4.17 19.88 4.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 17.95 3.5 19.4 3.8 ;
        RECT 19 3.45 19.3 3.8 ;
        RECT 19.05 1.85 19.3 3.8 ;
        RECT 17.95 1.85 19.3 2.1 ;
        RECT 17.95 3.5 18.2 5.2 ;
        RECT 17.95 0.95 18.2 2.1 ;
      LAYER MET2 ;
        RECT 18.9 3.5 19.4 3.8 ;
        RECT 18.95 3.45 19.35 3.85 ;
      LAYER VIA12 ;
        RECT 19.02 3.52 19.28 3.78 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.8 2.75 1.1 3.25 ;
      LAYER MET2 ;
        RECT 0.7 2.85 1.2 3.15 ;
        RECT 0.75 2.8 1.15 3.2 ;
      LAYER VIA12 ;
        RECT 0.82 2.87 1.08 3.13 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.9 2.85 16.4 3.15 ;
        RECT 3.4 3 3.9 3.3 ;
      LAYER MET2 ;
        RECT 15.9 2.8 16.4 3.2 ;
        RECT 3.5 4.95 16.3 5.25 ;
        RECT 16 2.8 16.3 5.25 ;
        RECT 3.4 2.95 3.9 3.35 ;
        RECT 3.5 2.95 3.8 5.25 ;
      LAYER VIA12 ;
        RECT 3.52 3.02 3.78 3.28 ;
        RECT 16.02 2.87 16.28 3.13 ;
    END
  END SN
  OBS
    LAYER MET2 ;
      RECT 18.15 2.5 18.55 2.9 ;
      RECT 18 2.55 18.6 2.85 ;
      RECT 16.6 2.05 16.9 2.55 ;
      RECT 2.65 2.15 3.15 2.55 ;
      RECT 1.35 2.15 1.75 2.55 ;
      RECT 16.55 2.05 16.95 2.5 ;
      RECT 1.3 2.2 3.15 2.5 ;
      RECT 2.75 0.9 3.05 2.55 ;
      RECT 16.55 0.9 16.85 2.5 ;
      RECT 2.75 0.9 16.85 1.2 ;
      RECT 10.7 1.5 11 4.05 ;
      RECT 10.65 3.6 11.05 4 ;
      RECT 14.6 2 15.1 2.4 ;
      RECT 14.6 1.55 15 2.4 ;
      RECT 10.65 1.5 11.05 1.9 ;
      RECT 10.6 1.55 15 1.85 ;
      RECT 12.4 4.15 12.8 4.55 ;
      RECT 12.35 4.2 14.5 4.5 ;
      RECT 14.2 2.85 14.5 4.5 ;
      RECT 12.45 2.4 12.75 4.55 ;
      RECT 14.2 2.85 15.05 3.2 ;
      RECT 14.55 2.8 15.05 3.2 ;
      RECT 12.4 2.4 12.8 2.8 ;
      RECT 12.35 2.45 12.85 2.75 ;
      RECT 7.1 4.35 11.7 4.65 ;
      RECT 11.4 2.15 11.7 4.65 ;
      RECT 7.1 2.1 7.4 4.65 ;
      RECT 11.35 2.2 11.75 2.6 ;
      RECT 7.05 2.1 7.5 2.5 ;
      RECT 7 2.15 7.5 2.45 ;
      RECT 9 1.5 9.3 2.4 ;
      RECT 8.95 1.95 9.35 2.35 ;
      RECT 8.95 2 9.4 2.3 ;
      RECT 4.65 1.85 5.15 2.25 ;
      RECT 4.65 1.9 6.6 2.2 ;
      RECT 6.3 1.5 6.6 2.2 ;
      RECT 8.95 1.5 9.3 2.35 ;
      RECT 6.3 1.5 9.3 1.8 ;
      RECT 4.4 2.95 4.9 3.35 ;
    LAYER VIA12 ;
      RECT 18.22 2.57 18.48 2.83 ;
      RECT 16.62 2.17 16.88 2.43 ;
      RECT 14.72 2.07 14.98 2.33 ;
      RECT 14.67 2.87 14.93 3.13 ;
      RECT 12.47 2.47 12.73 2.73 ;
      RECT 12.47 4.22 12.73 4.48 ;
      RECT 11.42 2.27 11.68 2.53 ;
      RECT 10.72 1.57 10.98 1.83 ;
      RECT 10.72 3.67 10.98 3.93 ;
      RECT 9.02 2.02 9.28 2.28 ;
      RECT 7.12 2.17 7.38 2.43 ;
      RECT 4.77 1.92 5.03 2.18 ;
      RECT 4.52 3.02 4.78 3.28 ;
      RECT 2.77 2.22 3.03 2.48 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 17.2 3.85 17.45 5.2 ;
      RECT 17.25 1.65 17.5 4.1 ;
      RECT 14.55 2.85 15.65 3.15 ;
      RECT 15.35 1.65 15.65 3.15 ;
      RECT 17.25 2.55 18.6 2.85 ;
      RECT 15.35 1.65 17.5 1.9 ;
      RECT 16.2 0.95 16.45 1.9 ;
      RECT 16.35 3.75 16.6 5.2 ;
      RECT 14.65 3.75 14.9 5.2 ;
      RECT 14.65 3.75 16.6 4 ;
      RECT 13.75 3.6 14 5.2 ;
      RECT 13.75 3.6 14.3 3.85 ;
      RECT 14.05 2.2 14.3 3.85 ;
      RECT 11.4 1.95 11.7 2.7 ;
      RECT 13.75 2.2 14.3 2.5 ;
      RECT 11.4 1.95 14 2.2 ;
      RECT 13.75 0.95 14 2.5 ;
      RECT 12.35 4.2 12.85 4.5 ;
      RECT 12.45 4.1 12.75 4.5 ;
      RECT 10.7 0.95 11 1.95 ;
      RECT 10.7 0.95 11.25 1.65 ;
      RECT 10.7 3.7 11.25 5.2 ;
      RECT 10.7 3.55 11 5.2 ;
      RECT 9 2 9.3 2.35 ;
      RECT 8.9 2 9.4 2.3 ;
      RECT 7.6 4.2 8.15 5.2 ;
      RECT 5.4 4.2 8.15 4.5 ;
      RECT 5.4 2.2 5.7 4.5 ;
      RECT 4.4 3 5.7 3.3 ;
      RECT 5.4 2.2 6.55 2.5 ;
      RECT 6.25 1.4 6.55 2.5 ;
      RECT 6.25 1.4 8.15 1.65 ;
      RECT 7.6 0.95 8.15 1.65 ;
      RECT 2.15 1.65 2.4 5.2 ;
      RECT 3.85 1.9 5.15 2.2 ;
      RECT 3.15 1.6 4.1 1.9 ;
      RECT 2.15 1.65 4.1 1.9 ;
      RECT 3.15 0.95 3.4 1.9 ;
      RECT 4.7 3.75 4.95 5.2 ;
      RECT 3 3.75 3.25 5.2 ;
      RECT 3 3.75 4.95 4 ;
      RECT 1.4 0.95 1.65 5.2 ;
      RECT 1.4 1.9 1.7 2.55 ;
      RECT 1.4 2.2 1.8 2.5 ;
      RECT 16.5 2.15 17 2.45 ;
      RECT 14.6 2.05 15.1 2.35 ;
      RECT 12.35 2.45 12.85 2.75 ;
      RECT 7 2.15 7.5 2.45 ;
      RECT 2.65 2.2 3.15 2.5 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffsr_1
