# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dff_1 0 0 ;
  SIZE 14.5 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 14.5 6.35 ;
        RECT 12.85 4.15 13.1 6.35 ;
        RECT 10.4 3.6 10.65 6.35 ;
        RECT 8.6 4.85 8.85 6.35 ;
        RECT 5 4.2 5.25 6.35 ;
        RECT 1.4 4.85 1.65 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 14.5 0.7 ;
        RECT 12.85 0 13.1 1.7 ;
        RECT 10.4 0 10.65 1.5 ;
        RECT 8.6 0 8.85 1.6 ;
        RECT 5 0 5.25 1.5 ;
        RECT 1.4 0 1.65 1.6 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 9 2.95 9.5 3.25 ;
        RECT 2.5 3.1 9.4 3.35 ;
        RECT 2.5 3.1 8.95 3.4 ;
        RECT 5.95 2.05 6.45 2.35 ;
        RECT 6.05 2.05 6.35 3.4 ;
        RECT 3.8 2.1 4.3 2.4 ;
        RECT 3.9 2.1 4.2 3.4 ;
      LAYER Metal2 ;
        RECT 9 2.95 9.5 3.25 ;
        RECT 9.05 2.9 9.45 3.3 ;
      LAYER Via1 ;
        RECT 9.12 2.97 9.38 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 2.95 2.25 3.25 ;
      LAYER Metal2 ;
        RECT 1.7 2.95 2.3 3.25 ;
        RECT 1.75 2.9 2.25 3.3 ;
      LAYER Via1 ;
        RECT 1.87 2.97 2.13 3.23 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.7 4.25 14.25 4.6 ;
        RECT 13.7 4.2 14.2 4.6 ;
        RECT 13.7 1.05 13.95 5.3 ;
      LAYER Metal2 ;
        RECT 13.75 4.25 14.25 4.55 ;
        RECT 13.8 4.2 14.2 4.6 ;
      LAYER Via1 ;
        RECT 13.87 4.27 14.13 4.53 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12 3.6 13.45 3.9 ;
        RECT 13.05 1.95 13.35 3.9 ;
        RECT 12 1.95 13.35 2.2 ;
        RECT 12 3.6 12.25 5.3 ;
        RECT 12 1.05 12.25 2.2 ;
      LAYER Metal2 ;
        RECT 12.95 3.6 13.45 3.9 ;
        RECT 13 3.55 13.4 3.95 ;
      LAYER Via1 ;
        RECT 13.07 3.62 13.33 3.88 ;
    END
  END QN
  OBS
    LAYER Metal2 ;
      RECT 8.1 4.25 8.5 4.65 ;
      RECT 8.05 4.3 11.45 4.6 ;
      RECT 11.15 2.65 11.45 4.6 ;
      RECT 8.15 2.25 8.45 4.65 ;
      RECT 12.2 2.6 12.6 3 ;
      RECT 11.15 2.65 12.65 2.95 ;
      RECT 8.1 2.25 8.5 2.65 ;
      RECT 8.05 2.3 8.55 2.6 ;
      RECT 6.5 1 6.8 4.7 ;
      RECT 6.45 4.25 6.85 4.65 ;
      RECT 10.55 1.7 10.95 2.1 ;
      RECT 10.2 1.75 11 2.05 ;
      RECT 6.45 1.4 6.85 1.8 ;
      RECT 6.5 1 6.85 1.8 ;
      RECT 10.2 1.7 10.95 2.05 ;
      RECT 10.2 1 10.5 2.05 ;
      RECT 6.5 1 10.5 1.3 ;
      RECT 2.8 5 7.55 5.3 ;
      RECT 7.25 1.6 7.55 5.3 ;
      RECT 2.8 2.05 3.1 5.3 ;
      RECT 2.75 2.05 3.2 2.45 ;
      RECT 2.7 2.1 3.2 2.4 ;
      RECT 9.4 1.6 9.8 2 ;
      RECT 7.2 1.6 7.6 2 ;
      RECT 7.15 1.65 9.9 1.95 ;
      RECT 4.65 2.05 5.05 2.45 ;
      RECT 0.45 2.05 0.85 2.45 ;
      RECT 4.6 2.1 5.1 2.4 ;
      RECT 0.4 2.1 0.9 2.4 ;
      RECT 4.7 1.15 5 2.45 ;
      RECT 0.5 1.15 0.8 2.45 ;
      RECT 0.5 1.15 5 1.45 ;
    LAYER Via1 ;
      RECT 12.27 2.67 12.53 2.93 ;
      RECT 10.62 1.77 10.88 2.03 ;
      RECT 9.47 1.67 9.73 1.93 ;
      RECT 8.17 2.32 8.43 2.58 ;
      RECT 8.17 4.32 8.43 4.58 ;
      RECT 7.27 1.67 7.53 1.93 ;
      RECT 6.52 1.47 6.78 1.73 ;
      RECT 6.52 4.32 6.78 4.58 ;
      RECT 4.72 2.12 4.98 2.38 ;
      RECT 2.82 2.12 3.08 2.38 ;
      RECT 0.52 2.12 0.78 2.38 ;
    LAYER Metal1 ;
      RECT 11.25 1.05 11.5 5.3 ;
      RECT 11.25 2.65 12.65 2.95 ;
      RECT 10.6 1.75 10.9 3.05 ;
      RECT 10.5 1.75 11 2.05 ;
      RECT 9.45 3.6 9.7 5.3 ;
      RECT 9.45 3.6 10 3.85 ;
      RECT 9.75 2.3 10 3.85 ;
      RECT 9.45 1.55 9.75 2.6 ;
      RECT 9.45 1.05 9.7 2.6 ;
      RECT 8.05 4.3 8.55 4.6 ;
      RECT 8.15 4.2 8.45 4.6 ;
      RECT 6.95 2 7.25 2.5 ;
      RECT 6.9 2.1 7.55 2.4 ;
      RECT 7.25 1.55 7.55 2.4 ;
      RECT 4.7 2.1 5 2.45 ;
      RECT 4.6 2.1 5.1 2.4 ;
      RECT 3.3 4.3 3.85 5.3 ;
      RECT 1.05 4.3 3.85 4.6 ;
      RECT 1.05 1.9 1.35 4.6 ;
      RECT 1.05 3.1 1.45 3.4 ;
      RECT 1.05 1.9 2.25 2.15 ;
      RECT 2 1.5 2.25 2.15 ;
      RECT 2 1.5 3.85 1.75 ;
      RECT 3.3 1.05 3.85 1.75 ;
      RECT 0.55 1.05 0.8 5.3 ;
      RECT 0.5 2 0.8 2.45 ;
      RECT 0.4 2.1 0.8 2.4 ;
      RECT 8.05 2.3 8.55 2.6 ;
      RECT 6.4 1.05 6.95 1.75 ;
      RECT 6.4 4.2 6.95 5.3 ;
      RECT 2.7 2.1 3.2 2.4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dff_1
