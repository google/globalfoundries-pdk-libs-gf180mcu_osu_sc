# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux2_1 0 0 ;
  SIZE 5.1 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 5.1 6.35 ;
        RECT 0.55 3.6 0.8 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.1 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 2.25 2.85 2.65 ;
        RECT 2.25 1.05 2.5 5.3 ;
      LAYER Metal2 ;
        RECT 2.35 2.25 2.85 2.65 ;
      LAYER Via1 ;
        RECT 2.47 2.32 2.73 2.58 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.25 2.25 4.75 2.65 ;
        RECT 4.25 1.05 4.5 5.3 ;
      LAYER Metal2 ;
        RECT 4.25 2.25 4.75 2.65 ;
      LAYER Via1 ;
        RECT 4.37 2.32 4.63 2.58 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 2.95 1.05 3.25 ;
      LAYER Metal2 ;
        RECT 0.55 2.9 1.05 3.3 ;
      LAYER Via1 ;
        RECT 0.67 2.97 0.93 3.23 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.1 4.15 3.4 4.65 ;
        RECT 3.1 1.05 3.35 5.3 ;
      LAYER Metal2 ;
        RECT 3 4.2 3.5 4.6 ;
      LAYER Via1 ;
        RECT 3.12 4.27 3.38 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 3.55 3.1 4.05 3.5 ;
      RECT 1.45 3.1 1.95 3.5 ;
      RECT 1.45 3.15 4.05 3.45 ;
    LAYER Via1 ;
      RECT 3.67 3.17 3.93 3.43 ;
      RECT 1.57 3.17 1.83 3.43 ;
    LAYER Metal1 ;
      RECT 1.4 1.05 1.65 5.3 ;
      RECT 1.4 3.15 1.95 3.45 ;
      RECT 1.4 2.1 2 2.4 ;
      RECT 3.65 3 3.95 3.55 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux2_1
