magic
tech gf180mcuC
timestamp 1661874610
<< error_p >>
rect 0 111 18 123
rect 2 61 18 111
rect 0 0 5 12
<< nwell >>
rect 0 61 2 123
<< metal1 >>
rect 0 111 2 123
rect 0 0 2 12
<< labels >>
rlabel metal1 1 117 1 117 3 VDD
rlabel metal1 1 5 1 5 2 GND
<< end >>
