* SKY130 Spice File.
.include "../../sky130_fd_pr__nfet_01v8__tt_leak.corner.spice"
.include "../../sky130_fd_pr__nfet_01v8__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_01v8_lvt__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__nfet_01v8_lvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__esd_nfet_01v8__tt_leak.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_lvt__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_lvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d10v5__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d10v5__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d10v5__mismatch.corner.spice"
.include "../../sky130_fd_pr__esd_pfet_g5v0d10v5__tt_leak.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_hvt__tt_leak.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8_hvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__pfet_01v8__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_05v0_nvt__tt_leak.corner.spice"
.include "../../sky130_fd_pr__nfet_05v0_nvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__nfet_g5v0d16v0__tt_leak_discrete.corner.spice"
.include "../../sky130_fd_pr__nfet_03v3_nvt__tt.corner.spice"
.include "../../sky130_fd_pr__nfet_03v3_nvt__mismatch.corner.spice"
.include "../../sky130_fd_pr__esd_nfet_g5v0d10v5__tt_leak.corner.spice"
.include "../../sky130_fd_pr__pfet_g5v0d16v0__tt_leak.corner.spice"
.include "nonfet.spice"
.include "../../all.spice"
.include "leakrf.spice"
