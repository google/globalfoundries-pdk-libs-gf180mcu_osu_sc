# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_nor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_nor2_1 0 0 ;
  SIZE 2.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.5 0.95 3.8 ;
      LAYER MET2 ;
        RECT 0.45 3.45 0.95 3.85 ;
      LAYER VIA12 ;
        RECT 0.57 3.52 0.83 3.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.85 2.85 2.35 3.15 ;
      LAYER MET2 ;
        RECT 1.85 2.8 2.35 3.2 ;
      LAYER VIA12 ;
        RECT 1.97 2.87 2.23 3.13 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
      LAYER MET2 ;
        RECT 1.65 7.55 2.15 7.85 ;
        RECT 1.7 7.5 2.1 7.9 ;
        RECT 0.45 7.55 0.95 7.85 ;
        RECT 0.5 7.5 0.9 7.9 ;
      LAYER VIA12 ;
        RECT 0.57 7.57 0.83 7.83 ;
        RECT 1.77 7.57 2.03 7.83 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 2.8 0.6 ;
        RECT 2.1 0 2.35 1.8 ;
        RECT 0.4 0 0.65 1.8 ;
      LAYER MET2 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 4.75 2.2 7.15 ;
        RECT 1.25 4.75 2.2 5 ;
        RECT 1.15 4.15 1.65 4.45 ;
        RECT 1.25 0.95 1.5 5 ;
      LAYER MET2 ;
        RECT 1.15 4.1 1.65 4.5 ;
      LAYER VIA12 ;
        RECT 1.27 4.17 1.53 4.43 ;
    END
  END Y
END gf180mcu_osu_sc_12T_nor2_1
