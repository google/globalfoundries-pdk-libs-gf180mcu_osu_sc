# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_xnor2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_xnor2_1 0 -0.15 ;
  SIZE 6.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.55 3.35 4.05 3.65 ;
        RECT 1.25 2.05 1.75 2.35 ;
      LAYER MET2 ;
        RECT 3.6 3.3 4 3.7 ;
        RECT 3.65 0.75 3.95 3.75 ;
        RECT 1.35 0.75 3.95 1.05 ;
        RECT 1.3 2 1.7 2.4 ;
        RECT 1.35 0.75 1.65 2.45 ;
      LAYER VIA12 ;
        RECT 1.37 2.07 1.63 2.33 ;
        RECT 3.67 3.37 3.93 3.63 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.35 2.05 4.85 2.35 ;
      LAYER MET2 ;
        RECT 4.35 2.05 4.85 2.35 ;
        RECT 4.4 2 4.8 2.4 ;
        RECT 4.45 1.95 4.75 2.45 ;
      LAYER VIA12 ;
        RECT 4.47 2.07 4.73 2.33 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 6.2 7.95 ;
        RECT 4.5 5.3 4.75 7.95 ;
        RECT 1.4 5.3 1.65 7.95 ;
      LAYER MET2 ;
        RECT 5.25 7.4 5.75 7.7 ;
        RECT 5.3 7.35 5.7 7.75 ;
        RECT 4.05 7.4 4.55 7.7 ;
        RECT 4.1 7.35 4.5 7.75 ;
        RECT 2.85 7.4 3.35 7.7 ;
        RECT 2.9 7.35 3.3 7.75 ;
        RECT 1.65 7.4 2.15 7.7 ;
        RECT 1.7 7.35 2.1 7.75 ;
        RECT 0.45 7.4 0.95 7.7 ;
        RECT 0.5 7.35 0.9 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
        RECT 1.77 7.42 2.03 7.68 ;
        RECT 2.97 7.42 3.23 7.68 ;
        RECT 4.17 7.42 4.43 7.68 ;
        RECT 5.37 7.42 5.63 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 6.2 0.45 ;
        RECT 4.5 -0.15 4.75 1.65 ;
        RECT 1.4 -0.15 1.65 1.65 ;
      LAYER MET2 ;
        RECT 5.25 0.1 5.75 0.4 ;
        RECT 5.3 0.05 5.7 0.45 ;
        RECT 4.05 0.1 4.55 0.4 ;
        RECT 4.1 0.05 4.5 0.45 ;
        RECT 2.85 0.1 3.35 0.4 ;
        RECT 2.9 0.05 3.3 0.45 ;
        RECT 1.65 0.1 2.15 0.4 ;
        RECT 1.7 0.05 2.1 0.45 ;
        RECT 0.45 0.1 0.95 0.4 ;
        RECT 0.5 0.05 0.9 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
        RECT 1.77 0.12 2.03 0.38 ;
        RECT 2.97 0.12 3.23 0.38 ;
        RECT 4.17 0.12 4.43 0.38 ;
        RECT 5.37 0.12 5.63 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 1.25 3.2 1.8 ;
        RECT 2.95 0.8 3.2 1.8 ;
        RECT 2.95 5.15 3.2 7 ;
        RECT 2.9 5.15 3.2 5.7 ;
      LAYER MET2 ;
        RECT 2.8 1.35 3.3 1.75 ;
        RECT 2.85 5.25 3.25 5.65 ;
        RECT 2.9 1.35 3.2 5.8 ;
      LAYER VIA12 ;
        RECT 2.92 5.32 3.18 5.58 ;
        RECT 2.92 1.42 3.18 1.68 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.35 0.8 5.6 7 ;
      RECT 2.55 4 5.6 4.3 ;
      RECT 0.55 0.8 0.8 7 ;
      RECT 0.55 3.35 3.3 3.65 ;
      RECT 3 2.05 3.3 3.65 ;
      RECT 2.9 2.05 3.4 2.35 ;
  END
END gf180mcu_osu_sc_12T_xnor2_1
