* NGSPICE file created from gf180mcu_osu_sc_12T_xnor2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y a_47_11# a_42_16# GND nmos_3p3 w=0.85u l=0.3u
X1 VDD B a_76_106# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_47_11# B VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 a_76_106# A Y VDD pmos_3p3 w=1.7u l=0.3u
X4 Y a_47_11# a_42_106# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_42_106# a_9_16# VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 VDD A a_9_16# VDD pmos_3p3 w=1.7u l=0.3u
X7 GND A a_9_16# GND nmos_3p3 w=0.85u l=0.3u
X8 a_76_16# a_9_16# Y GND nmos_3p3 w=0.85u l=0.3u
X9 a_42_16# A GND GND nmos_3p3 w=0.85u l=0.3u
X10 a_47_11# B GND GND nmos_3p3 w=0.85u l=0.3u
X11 GND B a_76_16# GND nmos_3p3 w=0.85u l=0.3u
