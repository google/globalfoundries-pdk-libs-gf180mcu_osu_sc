* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_aoi22_1 Y A0 A1 B0 B1
X0 a_9_109 B1 Y VDD pmos_3p3 w=34 l=6
X1 Y B0 a_9_109 VDD pmos_3p3 w=34 l=6
X2 a_9_109 A1 VDD VDD pmos_3p3 w=34 l=6
X3 VDD A0 a_9_109 VDD pmos_3p3 w=34 l=6
X4 a_56_19 B0 Y VSS nmos_3p3 w=17 l=6
X5 VSS B1 a_56_19 VSS nmos_3p3 w=17 l=6
X6 a_28_19 A0 VSS VSS nmos_3p3 w=17 l=6
X7 Y A1 a_28_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
