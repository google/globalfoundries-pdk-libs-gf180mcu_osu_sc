magic
tech gf180mcuC
timestamp 1660078683
<< nwell >>
rect 0 100 162 162
<< nmos >>
rect 19 19 25 36
rect 36 19 42 36
rect 53 19 59 36
rect 85 19 91 36
rect 102 19 108 36
rect 119 19 125 36
rect 136 19 142 36
<< pmos >>
rect 19 109 25 143
rect 36 109 42 143
rect 53 109 59 143
rect 85 109 91 143
rect 102 109 108 143
rect 119 109 125 143
rect 136 109 142 143
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 36 36
rect 25 21 28 34
rect 33 21 36 34
rect 25 19 36 21
rect 42 19 53 36
rect 59 34 69 36
rect 59 21 62 34
rect 67 21 69 34
rect 59 19 69 21
rect 75 34 85 36
rect 75 21 77 34
rect 82 21 85 34
rect 75 19 85 21
rect 91 34 102 36
rect 91 29 94 34
rect 99 29 102 34
rect 91 19 102 29
rect 108 34 119 36
rect 108 21 111 34
rect 116 21 119 34
rect 108 19 119 21
rect 125 34 136 36
rect 125 21 128 34
rect 133 21 136 34
rect 125 19 136 21
rect 142 34 152 36
rect 142 21 145 34
rect 150 21 152 34
rect 142 19 152 21
<< pdiff >>
rect 9 141 19 143
rect 9 111 11 141
rect 16 111 19 141
rect 9 109 19 111
rect 25 141 36 143
rect 25 111 28 141
rect 33 111 36 141
rect 25 109 36 111
rect 42 141 53 143
rect 42 111 45 141
rect 50 111 53 141
rect 42 109 53 111
rect 59 141 69 143
rect 59 111 62 141
rect 67 111 69 141
rect 59 109 69 111
rect 75 141 85 143
rect 75 111 77 141
rect 82 111 85 141
rect 75 109 85 111
rect 91 109 102 143
rect 108 141 119 143
rect 108 111 111 141
rect 116 111 119 141
rect 108 109 119 111
rect 125 141 136 143
rect 125 111 128 141
rect 133 111 136 141
rect 125 109 136 111
rect 142 141 152 143
rect 142 111 145 141
rect 150 111 152 141
rect 142 109 152 111
<< ndiffc >>
rect 11 21 16 34
rect 28 21 33 34
rect 62 21 67 34
rect 77 21 82 34
rect 94 29 99 34
rect 111 21 116 34
rect 128 21 133 34
rect 145 21 150 34
<< pdiffc >>
rect 11 111 16 141
rect 28 111 33 141
rect 45 111 50 141
rect 62 111 67 141
rect 77 111 82 141
rect 111 111 116 141
rect 128 111 133 141
rect 145 111 150 141
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
rect 81 10 90 12
rect 81 5 83 10
rect 88 5 90 10
rect 81 3 90 5
rect 105 10 114 12
rect 105 5 107 10
rect 112 5 114 10
rect 105 3 114 5
rect 129 10 138 12
rect 129 5 131 10
rect 136 5 138 10
rect 129 3 138 5
<< nsubdiff >>
rect 9 157 18 159
rect 9 152 11 157
rect 16 152 18 157
rect 9 150 18 152
rect 33 157 42 159
rect 33 152 35 157
rect 40 152 42 157
rect 33 150 42 152
rect 57 157 66 159
rect 57 152 59 157
rect 64 152 66 157
rect 57 150 66 152
rect 81 157 90 159
rect 81 152 83 157
rect 88 152 90 157
rect 81 150 90 152
rect 105 157 114 159
rect 105 152 107 157
rect 112 152 114 157
rect 105 150 114 152
rect 129 157 138 159
rect 129 152 131 157
rect 136 152 138 157
rect 129 150 138 152
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
rect 83 5 88 10
rect 107 5 112 10
rect 131 5 136 10
<< nsubdiffcont >>
rect 11 152 16 157
rect 35 152 40 157
rect 59 152 64 157
rect 83 152 88 157
rect 107 152 112 157
rect 131 152 136 157
<< polysilicon >>
rect 19 143 25 148
rect 36 143 42 148
rect 53 143 59 148
rect 85 143 91 148
rect 102 143 108 148
rect 119 143 125 148
rect 136 143 142 148
rect 19 104 25 109
rect 19 102 31 104
rect 19 96 23 102
rect 29 96 31 102
rect 19 94 31 96
rect 19 36 25 94
rect 36 78 42 109
rect 30 76 42 78
rect 30 70 32 76
rect 38 70 42 76
rect 30 68 42 70
rect 36 36 42 68
rect 53 65 59 109
rect 85 78 91 109
rect 78 76 91 78
rect 78 70 80 76
rect 86 70 91 76
rect 78 68 91 70
rect 47 63 59 65
rect 47 57 49 63
rect 55 57 59 63
rect 47 55 59 57
rect 53 36 59 55
rect 85 36 91 68
rect 102 65 108 109
rect 119 104 125 109
rect 119 102 131 104
rect 119 96 123 102
rect 129 96 131 102
rect 119 94 131 96
rect 102 63 114 65
rect 102 57 106 63
rect 112 57 114 63
rect 102 55 114 57
rect 102 36 108 55
rect 119 36 125 94
rect 136 78 142 109
rect 130 76 142 78
rect 130 70 132 76
rect 138 70 142 76
rect 130 68 142 70
rect 136 36 142 68
rect 19 14 25 19
rect 36 14 42 19
rect 53 14 59 19
rect 85 14 91 19
rect 102 14 108 19
rect 119 14 125 19
rect 136 14 142 19
<< polycontact >>
rect 23 96 29 102
rect 32 70 38 76
rect 80 70 86 76
rect 49 57 55 63
rect 123 96 129 102
rect 106 57 112 63
rect 132 70 138 76
<< metal1 >>
rect 0 157 162 162
rect 0 151 11 157
rect 17 151 35 157
rect 41 151 59 157
rect 65 151 83 157
rect 89 151 107 157
rect 113 151 131 157
rect 137 151 162 157
rect 0 150 162 151
rect 11 141 16 143
rect 11 50 16 111
rect 28 141 33 150
rect 28 109 33 111
rect 45 141 50 143
rect 45 102 50 111
rect 62 141 67 150
rect 62 109 67 111
rect 77 141 82 150
rect 77 109 82 111
rect 111 141 116 143
rect 21 96 23 102
rect 29 96 62 102
rect 68 96 70 102
rect 30 70 32 76
rect 38 70 40 76
rect 47 57 49 63
rect 55 57 57 63
rect 8 44 10 50
rect 16 44 18 50
rect 11 34 16 44
rect 11 19 16 21
rect 28 34 33 36
rect 28 12 33 21
rect 62 34 67 96
rect 111 76 116 111
rect 128 141 133 150
rect 128 109 133 111
rect 145 141 150 143
rect 145 103 150 111
rect 145 102 152 103
rect 121 96 123 102
rect 129 96 131 102
rect 144 96 146 102
rect 152 96 154 102
rect 145 95 152 96
rect 78 70 80 76
rect 86 70 88 76
rect 111 75 132 76
rect 94 70 132 75
rect 138 70 140 76
rect 62 19 67 21
rect 77 34 82 38
rect 94 34 99 70
rect 104 57 106 63
rect 112 57 114 63
rect 94 27 99 29
rect 111 34 116 38
rect 82 21 111 22
rect 77 17 116 21
rect 128 34 133 36
rect 128 12 133 21
rect 145 34 150 95
rect 145 19 150 21
rect 0 11 162 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 83 11
rect 89 5 107 11
rect 113 5 131 11
rect 137 5 162 11
rect 0 0 162 5
<< via1 >>
rect 11 152 16 157
rect 16 152 17 157
rect 11 151 17 152
rect 35 152 40 157
rect 40 152 41 157
rect 35 151 41 152
rect 59 152 64 157
rect 64 152 65 157
rect 59 151 65 152
rect 83 152 88 157
rect 88 152 89 157
rect 83 151 89 152
rect 107 152 112 157
rect 112 152 113 157
rect 107 151 113 152
rect 131 152 136 157
rect 136 152 137 157
rect 131 151 137 152
rect 62 96 68 102
rect 32 70 38 76
rect 49 57 55 63
rect 10 44 16 50
rect 123 96 129 102
rect 146 96 152 102
rect 80 70 86 76
rect 106 57 112 63
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
rect 83 10 89 11
rect 83 5 88 10
rect 88 5 89 10
rect 107 10 113 11
rect 107 5 112 10
rect 112 5 113 10
rect 131 10 137 11
rect 131 5 136 10
rect 136 5 137 10
<< metal2 >>
rect 10 157 18 158
rect 34 157 42 158
rect 58 157 66 158
rect 82 157 90 158
rect 106 157 114 158
rect 130 157 138 158
rect 9 151 11 157
rect 17 151 19 157
rect 33 151 35 157
rect 41 151 43 157
rect 57 151 59 157
rect 65 151 67 157
rect 81 151 83 157
rect 89 151 91 157
rect 105 151 107 157
rect 113 151 115 157
rect 129 151 131 157
rect 137 151 139 157
rect 10 150 18 151
rect 34 150 42 151
rect 58 150 66 151
rect 82 150 90 151
rect 106 150 114 151
rect 130 150 138 151
rect 60 102 70 103
rect 121 102 131 103
rect 60 96 62 102
rect 68 96 123 102
rect 129 96 131 102
rect 60 95 70 96
rect 121 95 131 96
rect 144 102 154 103
rect 144 96 146 102
rect 152 96 154 102
rect 144 95 154 96
rect 30 76 40 77
rect 78 76 88 77
rect 30 70 32 76
rect 38 70 80 76
rect 86 70 88 76
rect 30 69 40 70
rect 78 69 88 70
rect 47 63 57 64
rect 104 63 114 64
rect 47 57 49 63
rect 55 57 106 63
rect 112 57 114 63
rect 47 56 57 57
rect 104 56 114 57
rect 8 50 18 51
rect 8 44 10 50
rect 16 44 18 50
rect 8 43 18 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 81 5 83 11
rect 89 5 91 11
rect 105 5 107 11
rect 113 5 115 11
rect 129 5 131 11
rect 137 5 139 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
<< labels >>
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 14 154 14 154 1 VDD
rlabel metal2 12 47 12 47 1 CO
port 4 n
rlabel metal2 35 73 35 73 1 A
port 1 n
rlabel metal2 52 60 52 60 1 B
port 2 n
rlabel metal2 149 99 149 99 1 S
port 3 n
<< end >>
