* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_dff_1 D Q QN CLK
X0 a_42_70 D VDD VDD pmos_3p3 w=34 l=6
X1 a_125_19 a_53_38 a_114_70 VDD pmos_3p3 w=34 l=6
X2 a_86_70 a_53_38 a_19_14 VDD pmos_3p3 w=34 l=6
X3 VDD a_161_42 a_148_70 VDD pmos_3p3 w=34 l=6
X4 GND a_9_19 a_86_19 GND nmos_3p3 w=17 l=6
X5 a_19_14 a_53_38 a_42_19 GND nmos_3p3 w=17 l=6
X6 GND a_161_42 QN GND nmos_3p3 w=17 l=6
X7 VDD a_9_19 a_86_70 VDD pmos_3p3 w=34 l=6
X8 a_19_14 CLK a_42_70 VDD pmos_3p3 w=34 l=6
X9 VDD a_161_42 QN VDD pmos_3p3 w=34 l=6
X10 GND a_19_14 a_9_19 GND nmos_3p3 w=17 l=6
X11 a_53_38 CLK GND GND nmos_3p3 w=17 l=6
X12 VDD a_19_14 a_9_19 VDD pmos_3p3 w=34 l=6
X13 a_53_38 CLK VDD VDD pmos_3p3 w=34 l=6
X14 a_148_19 a_53_38 a_125_19 GND nmos_3p3 w=17 l=6
X15 Q QN GND GND nmos_3p3 w=17 l=6
X16 a_114_19 a_9_19 GND GND nmos_3p3 w=17 l=6
X17 a_161_42 a_125_19 GND GND nmos_3p3 w=17 l=6
X18 a_148_70 CLK a_125_19 VDD pmos_3p3 w=34 l=6
X19 Q QN VDD VDD pmos_3p3 w=34 l=6
X20 a_114_70 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X21 a_161_42 a_125_19 VDD VDD pmos_3p3 w=34 l=6
X22 a_42_19 D GND GND nmos_3p3 w=17 l=6
X23 a_125_19 CLK a_114_19 GND nmos_3p3 w=17 l=6
X24 a_86_19 CLK a_19_14 GND nmos_3p3 w=17 l=6
X25 GND a_161_42 a_148_19 GND nmos_3p3 w=17 l=6
.ends

