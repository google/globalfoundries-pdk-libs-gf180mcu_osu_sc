magic
tech gf180mcuC
timestamp 1659394494
<< nwell >>
rect 0 97 352 159
<< metal1 >>
rect 0 147 352 159
rect 0 -3 352 9
<< end >>
