* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp12t3v3__tinv_2 A Y EN EN_BAR
X0 a_36_19 A a_25_19 VSS nmos_3p3 w=17 l=6
X1 VSS a_36_19 Y VSS nmos_3p3 w=17 l=6
X2 a_36_19 A a_25_109 VDD pmos_3p3 w=34 l=6
X3 VSS a_36_19 a_36_19 VSS nmos_3p3 w=17 l=6
X4 a_25_109 EN_BAR VDD VDD pmos_3p3 w=34 l=6
X5 a_25_19 EN VSS VSS nmos_3p3 w=17 l=6
X6 Y a_36_19 VSS VSS nmos_3p3 w=17 l=6
X7 VDD a_36_19 Y VDD pmos_3p3 w=34 l=6
X8 Y a_36_19 VDD VDD pmos_3p3 w=34 l=6
X9 VDD a_36_19 a_36_19 VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
