* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__inv_8.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__inv_8 A Y VDD VSS
X0 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X1 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X2 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X3 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X4 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X5 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X8 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X9 Y A VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS A Y VSS nfet_03p3 w=0.85u l=0.3u
X13 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
X14 Y A VDD VDD pfet_03p3 w=1.7u l=0.3u
X15 VDD A Y VDD pfet_03p3 w=1.7u l=0.3u
.ends
