* NGSPICE file created from gf180mcu_osu_sc_12T_dffn_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 a_19_11# CLKN a_42_106# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_75_106# a_52_11# a_19_11# VDD pmos_3p3 w=1.7u l=0.3u
X2 a_135_65# a_114_16# VDD VDD pmos_3p3 w=1.7u l=0.3u
X3 Q QN GND GND nmos_3p3 w=0.85u l=0.3u
X4 a_131_16# a_52_11# a_114_16# GND nmos_3p3 w=0.85u l=0.3u
X5 a_42_106# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X6 a_135_65# a_114_16# GND GND nmos_3p3 w=0.85u l=0.3u
X7 VDD a_19_11# a_9_16# VDD pmos_3p3 w=1.7u l=0.3u
X8 a_75_16# CLKN a_19_11# GND nmos_3p3 w=0.85u l=0.3u
X9 GND a_135_65# a_131_16# GND nmos_3p3 w=0.85u l=0.3u
X10 a_19_11# a_52_11# a_42_16# GND nmos_3p3 w=0.85u l=0.3u
X11 GND a_19_11# a_9_16# GND nmos_3p3 w=0.85u l=0.3u
X12 a_52_11# CLKN VDD VDD pmos_3p3 w=1.7u l=0.3u
X13 VDD a_135_65# a_131_106# VDD pmos_3p3 w=1.7u l=0.3u
X14 a_131_106# CLKN a_114_16# VDD pmos_3p3 w=1.7u l=0.3u
X15 GND a_135_65# QN GND nmos_3p3 w=0.85u l=0.3u
X16 a_114_16# a_52_11# a_103_106# VDD pmos_3p3 w=1.7u l=0.3u
X17 a_114_16# CLKN a_103_16# GND nmos_3p3 w=0.85u l=0.3u
X18 a_52_11# CLKN GND GND nmos_3p3 w=0.85u l=0.3u
X19 a_42_16# D GND GND nmos_3p3 w=0.85u l=0.3u
X20 VDD a_9_16# a_75_106# VDD pmos_3p3 w=1.7u l=0.3u
X21 a_103_106# a_9_16# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 a_103_16# a_9_16# GND GND nmos_3p3 w=0.85u l=0.3u
X23 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X24 VDD a_135_65# QN VDD pmos_3p3 w=1.7u l=0.3u
X25 GND a_9_16# a_75_16# GND nmos_3p3 w=0.85u l=0.3u
