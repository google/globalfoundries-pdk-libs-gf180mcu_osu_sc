* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_addh_1 A B S CO
X0 VDD B a_19_14 VDD pmos_3p3 w=34 l=6
X1 a_19_14 A VDD VDD pmos_3p3 w=34 l=6
X2 VDD a_19_14 CO VDD pmos_3p3 w=34 l=6
X3 a_19_14 B a_42_19 VSS nmos_3p3 w=17 l=6
X4 S a_91_19 VSS VSS nmos_3p3 w=17 l=6
X5 VSS a_19_14 CO VSS nmos_3p3 w=17 l=6
X6 S a_91_19 VDD VDD pmos_3p3 w=34 l=6
X7 a_91_19 B a_91_109 VDD pmos_3p3 w=34 l=6
X8 VDD a_19_14 a_91_19 VDD pmos_3p3 w=34 l=6
X9 a_91_109 A VDD VDD pmos_3p3 w=34 l=6
X10 a_91_19 A a_75_19 VSS nmos_3p3 w=17 l=6
X11 a_42_19 A VSS VSS nmos_3p3 w=17 l=6
X12 VSS a_19_14 a_75_19 VSS nmos_3p3 w=17 l=6
X13 a_75_19 B a_91_19 VSS nmos_3p3 w=17 l=6
.ends

** hspice subcircuit dictionary
