magic
tech gf180mcuC
timestamp 1661874504
<< nwell >>
rect 0 61 64 123
<< nmos >>
rect 19 19 25 36
rect 38 19 44 36
<< pmos >>
rect 19 70 25 104
rect 38 70 44 104
<< ndiff >>
rect 9 34 19 36
rect 9 21 11 34
rect 16 21 19 34
rect 9 19 19 21
rect 25 34 38 36
rect 25 21 28 34
rect 35 21 38 34
rect 25 19 38 21
rect 44 34 54 36
rect 44 21 47 34
rect 52 21 54 34
rect 44 19 54 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 102 38 104
rect 25 72 28 102
rect 35 72 38 102
rect 25 70 38 72
rect 44 102 54 104
rect 44 88 47 102
rect 52 88 54 102
rect 44 70 54 88
<< ndiffc >>
rect 11 21 16 34
rect 28 21 35 34
rect 47 21 52 34
<< pdiffc >>
rect 11 72 16 102
rect 28 72 35 102
rect 47 88 52 102
<< psubdiff >>
rect 9 10 19 12
rect 9 5 11 10
rect 16 5 19 10
rect 9 3 19 5
rect 33 10 43 12
rect 33 5 35 10
rect 40 5 43 10
rect 33 3 43 5
<< nsubdiff >>
rect 9 118 19 120
rect 9 113 11 118
rect 16 113 19 118
rect 9 111 19 113
rect 33 118 43 120
rect 33 113 35 118
rect 40 113 43 118
rect 33 111 43 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
<< polysilicon >>
rect 19 104 25 109
rect 38 104 44 109
rect 19 65 25 70
rect 19 63 31 65
rect 19 57 23 63
rect 29 57 31 63
rect 19 55 31 57
rect 19 36 25 55
rect 38 51 44 70
rect 34 49 44 51
rect 34 43 36 49
rect 42 43 44 49
rect 34 41 44 43
rect 38 36 44 41
rect 19 14 25 19
rect 38 14 44 19
<< polycontact >>
rect 23 57 29 63
rect 36 43 42 49
<< metal1 >>
rect 0 118 64 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 64 118
rect 0 111 64 112
rect 11 102 16 104
rect 11 49 16 72
rect 28 102 35 111
rect 47 102 52 104
rect 47 76 52 88
rect 28 70 35 72
rect 45 70 47 76
rect 53 70 55 76
rect 21 57 23 63
rect 29 57 31 63
rect 11 43 36 49
rect 42 43 44 49
rect 11 34 16 43
rect 11 19 16 21
rect 28 34 35 36
rect 45 30 47 36
rect 53 30 55 36
rect 28 12 35 21
rect 47 19 52 21
rect 0 11 64 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 64 11
rect 0 0 64 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 47 70 53 76
rect 23 57 29 63
rect 47 34 53 36
rect 47 30 52 34
rect 52 30 53 34
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 10 111 18 112
rect 34 111 42 112
rect 45 76 55 77
rect 45 70 47 76
rect 53 70 55 76
rect 45 69 55 70
rect 22 63 30 64
rect 21 57 23 63
rect 29 57 31 63
rect 22 56 30 57
rect 47 37 53 69
rect 45 36 55 37
rect 45 30 47 36
rect 53 30 55 36
rect 45 29 55 30
rect 10 11 18 12
rect 34 11 42 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 10 4 18 5
rect 34 4 42 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 26 60 26 60 1 A
port 1 n
rlabel metal2 50 73 50 73 1 Y
port 2 n
<< end >>
