# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__lshifdown
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifdown 0 0 ;
  SIZE 5.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 7.6 5.2 8.3 ;
        RECT 3.45 5.55 3.75 8.3 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.3 8.3 ;
        RECT 0.55 5.55 0.85 8.3 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.2 0.7 ;
        RECT 3.45 0 3.75 1.9 ;
        RECT 0.55 0 0.85 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.3 4.25 4.7 4.55 ;
        RECT 4.35 1.05 4.65 7.25 ;
      LAYER Metal2 ;
        RECT 4.25 4.2 4.75 4.6 ;
      LAYER Via1 ;
        RECT 4.37 4.27 4.63 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 3.5 4.85 4 5.25 ;
      RECT 1.35 4.85 1.85 5.25 ;
      RECT 1.35 4.9 4 5.2 ;
    LAYER Via1 ;
      RECT 3.62 4.92 3.88 5.18 ;
      RECT 1.47 4.92 1.73 5.18 ;
    LAYER Metal1 ;
      RECT 1.45 1.05 1.75 7.25 ;
      RECT 1.35 4.9 1.85 5.2 ;
      RECT 3.5 4.9 4 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifdown
