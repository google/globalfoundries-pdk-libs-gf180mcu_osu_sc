# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__aoi22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi22_1 0 0 ;
  SIZE 5.35 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.35 8.3 ;
        RECT 1.4 6.3 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.35 0.7 ;
        RECT 3.5 0 3.75 1.9 ;
        RECT 0.7 0 0.95 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 3.6 1.1 3.9 ;
      LAYER Metal2 ;
        RECT 0.6 3.55 1.1 3.95 ;
      LAYER Via1 ;
        RECT 0.72 3.62 0.98 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 4.25 2.1 4.55 ;
      LAYER Metal2 ;
        RECT 1.6 4.2 2.1 4.6 ;
      LAYER Via1 ;
        RECT 1.72 4.27 1.98 4.53 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.35 3.6 2.85 3.9 ;
      LAYER Metal2 ;
        RECT 2.35 3.55 2.85 3.95 ;
      LAYER Via1 ;
        RECT 2.47 3.62 2.73 3.88 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.3 4.25 3.8 4.55 ;
      LAYER Metal2 ;
        RECT 3.3 4.2 3.8 4.6 ;
      LAYER Via1 ;
        RECT 3.42 4.27 3.68 4.53 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.3 4.9 4.8 5.2 ;
        RECT 4.45 6.1 4.75 6.6 ;
        RECT 4.45 4.9 4.7 6.6 ;
        RECT 4.4 3.1 4.65 5.2 ;
        RECT 2.1 3.1 4.65 3.35 ;
        RECT 2.1 1.05 2.35 3.35 ;
        RECT 3 6.2 3.5 6.5 ;
        RECT 3.1 6.2 3.35 7.25 ;
      LAYER Metal2 ;
        RECT 4.35 6.15 4.85 6.55 ;
        RECT 3 6.2 4.85 6.5 ;
        RECT 3 6.15 3.5 6.55 ;
        RECT 4.3 4.85 4.8 5.25 ;
      LAYER Via1 ;
        RECT 3.12 6.22 3.38 6.48 ;
        RECT 4.42 4.92 4.68 5.18 ;
        RECT 4.47 6.22 4.73 6.48 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 3.95 5.7 4.2 7.25 ;
      RECT 2.25 5.7 2.5 7.25 ;
      RECT 0.55 5.7 0.8 7.25 ;
      RECT 0.55 5.7 4.2 5.95 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi22_1
