* NGSPICE file created from gf180mcu_osu_sc_12T_tiehi.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y a_19_11# VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_11# a_19_11# GND GND nmos_3p3 w=0.85u l=0.3u
