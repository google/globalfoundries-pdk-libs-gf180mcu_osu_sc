magic
tech gf180mcuC
timestamp 1660079235
<< error_p >>
rect 0 147 18 159
rect 4 97 18 147
rect 0 -3 5 9
<< nwell >>
rect 0 97 4 159
<< metal1 >>
rect 0 147 4 159
rect 0 -3 4 9
<< labels >>
rlabel metal1 2 2 2 2 2 GND
rlabel metal1 2 152 2 152 3 VDD
<< end >>
