# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai21_1 0 0 ;
  SIZE 3.9 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 3.9 8.3 ;
        RECT 2.95 5.55 3.2 8.3 ;
        RECT 0.65 5.55 0.9 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.9 0.7 ;
        RECT 1.35 0 1.6 1.6 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.45 3.6 0.95 3.9 ;
      LAYER Metal2 ;
        RECT 0.45 3.55 0.95 3.95 ;
      LAYER Via1 ;
        RECT 0.57 3.62 0.83 3.88 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.45 4.25 1.95 4.55 ;
      LAYER Metal2 ;
        RECT 1.45 4.2 1.95 4.6 ;
      LAYER Via1 ;
        RECT 1.57 4.27 1.83 4.53 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.2 3.6 2.7 3.9 ;
      LAYER Metal2 ;
        RECT 2.2 3.55 2.7 3.95 ;
      LAYER Via1 ;
        RECT 2.32 3.62 2.58 3.88 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 4.9 3.35 5.2 ;
        RECT 3.05 1.05 3.3 2.6 ;
        RECT 2.95 2.35 3.2 5.2 ;
        RECT 2.1 4.9 2.35 7.25 ;
      LAYER Metal2 ;
        RECT 2.85 4.85 3.35 5.25 ;
      LAYER Via1 ;
        RECT 2.97 4.92 3.23 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.5 1.85 2.45 2.1 ;
      RECT 2.2 1.05 2.45 2.1 ;
      RECT 0.5 1.05 0.75 2.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai21_1
