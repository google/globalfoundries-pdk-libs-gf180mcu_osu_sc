# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_addf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_addf_1 0 0 ;
  SIZE 14 BY 6.15 ;
  SYMMETRY X Y ;
  SITE 9T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 8.7 2.35 9.2 2.65 ;
        RECT 6.4 3.05 9.1 3.35 ;
        RECT 8.8 2.35 9.1 3.35 ;
        RECT 6.4 2.35 6.7 3.35 ;
        RECT 3.2 2.35 6.7 2.65 ;
        RECT 2.15 3.1 3.45 3.4 ;
        RECT 3.2 2.35 3.45 3.4 ;
        RECT 2.15 2.2 2.4 3.4 ;
        RECT 0.6 2.2 2.4 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.85 3.6 9.95 3.9 ;
        RECT 9.65 2.9 9.95 3.9 ;
        RECT 5.85 2.9 6.15 3.9 ;
        RECT 3.7 3 6.15 3.3 ;
        RECT 1.6 3.65 4 3.95 ;
        RECT 3.7 2.9 4 3.95 ;
        RECT 1.6 2.75 1.9 3.95 ;
      LAYER MET2 ;
        RECT 1.5 2.85 2 3.15 ;
        RECT 1.55 2.8 1.95 3.2 ;
      LAYER VIA12 ;
        RECT 1.62 2.87 1.88 3.13 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 9.75 2.25 10.6 2.55 ;
        RECT 9.75 1.8 10.05 2.55 ;
        RECT 2.65 1.8 10.05 2.1 ;
        RECT 7.05 1.8 7.35 2.75 ;
        RECT 2.65 1.8 2.95 2.6 ;
      LAYER MET2 ;
        RECT 2.55 2.2 3.05 2.5 ;
        RECT 2.6 2.15 3 2.55 ;
      LAYER VIA12 ;
        RECT 2.67 2.22 2.93 2.48 ;
    END
  END CI
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.2 3 13.75 3.3 ;
        RECT 13.2 2.95 13.65 3.35 ;
        RECT 13.2 0.95 13.45 5.2 ;
      LAYER MET2 ;
        RECT 13.25 3 13.75 3.3 ;
        RECT 13.3 2.95 13.7 3.35 ;
      LAYER VIA12 ;
        RECT 13.37 3.02 13.63 3.28 ;
    END
  END CO
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14 0.6 ;
        RECT 12.35 0 12.6 1.4 ;
        RECT 10.75 0 11 1.4 ;
        RECT 6.5 0 6.75 1.4 ;
        RECT 4.8 0 5.05 1.4 ;
        RECT 1.4 0 1.65 1.4 ;
      LAYER MET2 ;
        RECT 12.45 0.25 12.95 0.55 ;
        RECT 12.5 0.2 12.9 0.6 ;
        RECT 11.25 0.25 11.75 0.55 ;
        RECT 11.3 0.2 11.7 0.6 ;
        RECT 10.05 0.25 10.55 0.55 ;
        RECT 10.1 0.2 10.5 0.6 ;
        RECT 8.85 0.25 9.35 0.55 ;
        RECT 8.9 0.2 9.3 0.6 ;
        RECT 7.65 0.25 8.15 0.55 ;
        RECT 7.7 0.2 8.1 0.6 ;
        RECT 6.45 0.25 6.95 0.55 ;
        RECT 6.5 0.2 6.9 0.6 ;
        RECT 5.25 0.25 5.75 0.55 ;
        RECT 5.3 0.2 5.7 0.6 ;
        RECT 4.05 0.25 4.55 0.55 ;
        RECT 4.1 0.2 4.5 0.6 ;
        RECT 2.85 0.25 3.35 0.55 ;
        RECT 2.9 0.2 3.3 0.6 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
        RECT 2.97 0.27 3.23 0.53 ;
        RECT 4.17 0.27 4.43 0.53 ;
        RECT 5.37 0.27 5.63 0.53 ;
        RECT 6.57 0.27 6.83 0.53 ;
        RECT 7.77 0.27 8.03 0.53 ;
        RECT 8.97 0.27 9.23 0.53 ;
        RECT 10.17 0.27 10.43 0.53 ;
        RECT 11.37 0.27 11.63 0.53 ;
        RECT 12.57 0.27 12.83 0.53 ;
    END
  END GND
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 11.6 3 12.05 3.3 ;
        RECT 11.6 2.95 11.9 3.35 ;
        RECT 11.6 0.95 11.85 5.2 ;
      LAYER MET2 ;
        RECT 11.55 3 12.05 3.3 ;
        RECT 11.6 2.95 12 3.35 ;
      LAYER VIA12 ;
        RECT 11.67 3.02 11.93 3.28 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 14 6.15 ;
        RECT 12.35 4.7 12.6 6.15 ;
        RECT 10.75 4.7 11 6.15 ;
        RECT 6.5 4.7 6.75 6.15 ;
        RECT 4.8 4.7 5.05 6.15 ;
        RECT 1.4 4.7 1.65 6.15 ;
      LAYER MET2 ;
        RECT 12.45 5.6 12.95 5.9 ;
        RECT 12.5 5.55 12.9 5.95 ;
        RECT 11.25 5.6 11.75 5.9 ;
        RECT 11.3 5.55 11.7 5.95 ;
        RECT 10.05 5.6 10.55 5.9 ;
        RECT 10.1 5.55 10.5 5.95 ;
        RECT 8.85 5.6 9.35 5.9 ;
        RECT 8.9 5.55 9.3 5.95 ;
        RECT 7.65 5.6 8.15 5.9 ;
        RECT 7.7 5.55 8.1 5.95 ;
        RECT 6.45 5.6 6.95 5.9 ;
        RECT 6.5 5.55 6.9 5.95 ;
        RECT 5.25 5.6 5.75 5.9 ;
        RECT 5.3 5.55 5.7 5.95 ;
        RECT 4.05 5.6 4.55 5.9 ;
        RECT 4.1 5.55 4.5 5.95 ;
        RECT 2.85 5.6 3.35 5.9 ;
        RECT 2.9 5.55 3.3 5.95 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
        RECT 2.97 5.62 3.23 5.88 ;
        RECT 4.17 5.62 4.43 5.88 ;
        RECT 5.37 5.62 5.63 5.88 ;
        RECT 6.57 5.62 6.83 5.88 ;
        RECT 7.77 5.62 8.03 5.88 ;
        RECT 8.97 5.62 9.23 5.88 ;
        RECT 10.17 5.62 10.43 5.88 ;
        RECT 11.37 5.62 11.63 5.88 ;
        RECT 12.57 5.62 12.83 5.88 ;
    END
  END VDD
  OBS
    LAYER MET2 ;
      RECT 3.1 4.75 3.4 5.2 ;
      RECT 3.05 4.75 3.45 5.15 ;
      RECT 3 4.8 12.85 5.1 ;
      RECT 12.55 2.25 12.85 5.1 ;
      RECT 3.75 1.05 4.05 5.1 ;
      RECT 12.5 2.3 12.9 2.7 ;
      RECT 7.85 2.3 8.25 2.7 ;
      RECT 12.45 2.35 12.95 2.65 ;
      RECT 3.75 2.35 8.3 2.65 ;
      RECT 3.1 0.95 3.4 1.45 ;
      RECT 3.05 1 3.45 1.4 ;
      RECT 3.05 1.05 4.05 1.35 ;
      RECT 8.15 4.1 8.55 4.5 ;
      RECT 8.1 4.15 11.25 4.45 ;
      RECT 10.95 2.25 11.25 4.45 ;
      RECT 8.85 1.05 9.15 4.45 ;
      RECT 10.9 2.3 11.3 2.7 ;
      RECT 8.15 1 8.55 1.4 ;
      RECT 8.1 1.05 9.15 1.35 ;
      RECT 7.3 0.95 7.6 1.45 ;
      RECT 5.65 0.95 5.95 1.45 ;
      RECT 7.25 1 7.65 1.4 ;
      RECT 5.6 1 6 1.4 ;
      RECT 5.6 1.05 7.65 1.35 ;
      RECT 2.2 0.95 2.5 1.45 ;
      RECT 0.5 0.95 0.8 1.45 ;
      RECT 2.15 1 2.55 1.4 ;
      RECT 0.45 1 0.85 1.4 ;
      RECT 0.45 1.05 2.55 1.35 ;
    LAYER VIA12 ;
      RECT 12.57 2.37 12.83 2.63 ;
      RECT 10.97 2.37 11.23 2.63 ;
      RECT 8.22 1.07 8.48 1.33 ;
      RECT 8.22 4.17 8.48 4.43 ;
      RECT 7.92 2.37 8.18 2.63 ;
      RECT 7.32 1.07 7.58 1.33 ;
      RECT 5.67 1.07 5.93 1.33 ;
      RECT 3.12 1.07 3.38 1.33 ;
      RECT 3.12 4.82 3.38 5.08 ;
      RECT 2.22 1.07 2.48 1.33 ;
      RECT 0.52 1.07 0.78 1.33 ;
    LAYER MET1 ;
      RECT 7.35 4.2 7.6 5.2 ;
      RECT 5.65 4.2 5.9 5.2 ;
      RECT 5.65 4.2 7.6 4.45 ;
      RECT 2.25 4.2 2.5 5.2 ;
      RECT 0.55 4.2 0.8 5.2 ;
      RECT 0.55 4.2 2.5 4.45 ;
      RECT 12.45 2.35 12.95 2.65 ;
      RECT 10.85 2.35 11.35 2.65 ;
      RECT 8.1 4.15 8.6 4.45 ;
      RECT 8.2 0.95 8.5 1.45 ;
      RECT 7.8 2.35 8.3 2.65 ;
      RECT 7.3 0.95 7.6 1.45 ;
      RECT 5.65 0.95 5.95 1.45 ;
      RECT 3.1 0.95 3.4 1.45 ;
      RECT 3.1 4.7 3.4 5.2 ;
      RECT 2.2 0.95 2.5 1.45 ;
      RECT 0.5 0.95 0.8 1.45 ;
  END
END gf180mcu_osu_sc_9T_addf_1
