// Copyright 2022 Google LLC
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
`timescale 1ns/10ps
`celldefine
module gf180mcu_osu_sc_9T_oai22_1 (Y, A0, A1);
	output Y;
	input A0, A1;

	// Function
	wire A0__bar, A1__bar;

	not (A1__bar, A1);
	not (A0__bar, A0);
	and (Y, A0__bar, A1__bar);

	// Timing
	specify
		(A0 => Y) = 0;
		(A1 => Y) = 0;
	endspecify
endmodule
`endcelldefine
