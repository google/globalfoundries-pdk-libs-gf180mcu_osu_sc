# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dffsr_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dffsr_1 0 0 ;
  SIZE 20.5 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 20.5 6.35 ;
        RECT 18.8 4.15 19.05 6.35 ;
        RECT 15.5 4.35 15.75 6.35 ;
        RECT 12.9 4.85 13.15 6.35 ;
        RECT 9.3 4.2 9.55 6.35 ;
        RECT 5.7 4.85 5.95 6.35 ;
        RECT 3.85 4.35 4.1 6.35 ;
        RECT 0.55 3.6 0.8 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 20.5 0.7 ;
        RECT 18.8 0 19.05 1.7 ;
        RECT 17.05 0 17.3 1.5 ;
        RECT 14.8 0 15.05 1.9 ;
        RECT 12.9 0 13.15 1.8 ;
        RECT 9.3 0 9.55 1.5 ;
        RECT 5.7 0 5.95 1.6 ;
        RECT 4.55 0 4.8 1.55 ;
        RECT 2.3 0 2.55 1.5 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 13.3 2.95 13.8 3.25 ;
        RECT 6.8 3.1 13.7 3.4 ;
        RECT 10.25 2.3 10.75 2.55 ;
        RECT 10.35 2.3 10.65 3.4 ;
        RECT 8.1 2.25 8.6 2.55 ;
        RECT 8.2 2.25 8.5 3.4 ;
      LAYER Metal2 ;
        RECT 13.3 2.95 13.8 3.25 ;
        RECT 13.35 2.9 13.75 3.3 ;
      LAYER Via1 ;
        RECT 13.42 2.97 13.68 3.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.05 2.95 6.55 3.25 ;
      LAYER Metal2 ;
        RECT 6 2.95 6.6 3.25 ;
        RECT 6.05 2.9 6.55 3.3 ;
      LAYER Via1 ;
        RECT 6.17 2.97 6.43 3.23 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 19.65 1.05 19.9 5.3 ;
        RECT 19.6 4.15 19.9 4.65 ;
      LAYER Metal2 ;
        RECT 19.5 4.25 20 4.55 ;
        RECT 19.55 4.2 19.95 4.6 ;
      LAYER Via1 ;
        RECT 19.62 4.27 19.88 4.53 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 17.95 3.6 19.4 3.9 ;
        RECT 19 3.55 19.3 3.9 ;
        RECT 19.05 1.95 19.3 3.9 ;
        RECT 17.95 1.95 19.3 2.2 ;
        RECT 17.95 3.6 18.2 5.3 ;
        RECT 17.95 1.05 18.2 2.2 ;
      LAYER Metal2 ;
        RECT 18.9 3.6 19.4 3.9 ;
        RECT 18.95 3.55 19.35 3.95 ;
      LAYER Via1 ;
        RECT 19.02 3.62 19.28 3.88 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 2.85 1.1 3.35 ;
      LAYER Metal2 ;
        RECT 0.7 2.95 1.2 3.25 ;
        RECT 0.75 2.9 1.15 3.3 ;
      LAYER Via1 ;
        RECT 0.82 2.97 1.08 3.23 ;
    END
  END RN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15.9 2.95 16.4 3.25 ;
        RECT 3.4 3.1 3.9 3.4 ;
      LAYER Metal2 ;
        RECT 15.9 2.9 16.4 3.3 ;
        RECT 3.5 5.05 16.3 5.35 ;
        RECT 16 2.9 16.3 5.35 ;
        RECT 3.4 3.05 3.9 3.45 ;
        RECT 3.5 3.05 3.8 5.35 ;
      LAYER Via1 ;
        RECT 3.52 3.12 3.78 3.38 ;
        RECT 16.02 2.97 16.28 3.23 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 18.15 2.6 18.55 3 ;
      RECT 18 2.65 18.6 2.95 ;
      RECT 16.6 2.15 16.9 2.65 ;
      RECT 2.65 2.25 3.15 2.65 ;
      RECT 1.35 2.25 1.75 2.65 ;
      RECT 16.55 2.15 16.95 2.6 ;
      RECT 1.3 2.3 3.15 2.6 ;
      RECT 2.75 1 3.05 2.65 ;
      RECT 16.55 1 16.85 2.6 ;
      RECT 2.75 1 16.85 1.3 ;
      RECT 10.8 1.6 11.1 4.15 ;
      RECT 10.75 3.7 11.15 4.1 ;
      RECT 14.6 2.1 15.1 2.5 ;
      RECT 14.6 1.65 15 2.5 ;
      RECT 10.75 1.6 11.15 2 ;
      RECT 10.7 1.65 15 1.95 ;
      RECT 12.4 4.25 12.8 4.65 ;
      RECT 12.35 4.3 14.5 4.6 ;
      RECT 14.2 2.95 14.5 4.6 ;
      RECT 12.45 2.5 12.75 4.65 ;
      RECT 14.2 2.95 15.05 3.3 ;
      RECT 14.55 2.9 15.05 3.3 ;
      RECT 12.4 2.5 12.8 2.9 ;
      RECT 12.35 2.55 12.85 2.85 ;
      RECT 7.1 4.45 11.8 4.75 ;
      RECT 11.5 2.25 11.8 4.75 ;
      RECT 7.1 2.2 7.4 4.75 ;
      RECT 11.45 2.3 11.85 2.7 ;
      RECT 7.05 2.2 7.5 2.6 ;
      RECT 7 2.25 7.5 2.55 ;
      RECT 9 1.6 9.3 2.5 ;
      RECT 8.95 2.05 9.35 2.45 ;
      RECT 8.95 2.1 9.4 2.4 ;
      RECT 4.65 1.95 5.15 2.35 ;
      RECT 4.65 2 6.6 2.3 ;
      RECT 6.3 1.6 6.6 2.3 ;
      RECT 8.95 1.6 9.3 2.45 ;
      RECT 6.3 1.6 9.3 1.9 ;
      RECT 4.4 3.05 4.9 3.45 ;
    LAYER Via1 ;
      RECT 18.22 2.67 18.48 2.93 ;
      RECT 16.62 2.27 16.88 2.53 ;
      RECT 14.72 2.17 14.98 2.43 ;
      RECT 14.67 2.97 14.93 3.23 ;
      RECT 12.47 2.57 12.73 2.83 ;
      RECT 12.47 4.32 12.73 4.58 ;
      RECT 11.52 2.37 11.78 2.63 ;
      RECT 10.82 1.67 11.08 1.93 ;
      RECT 10.82 3.77 11.08 4.03 ;
      RECT 9.02 2.12 9.28 2.38 ;
      RECT 7.12 2.27 7.38 2.53 ;
      RECT 4.77 2.02 5.03 2.28 ;
      RECT 4.52 3.12 4.78 3.38 ;
      RECT 2.77 2.32 3.03 2.58 ;
      RECT 1.42 2.32 1.68 2.58 ;
    LAYER Metal1 ;
      RECT 17.2 3.95 17.45 5.3 ;
      RECT 17.25 1.75 17.5 4.2 ;
      RECT 14.55 2.95 15.65 3.25 ;
      RECT 15.35 1.75 15.65 3.25 ;
      RECT 17.25 2.65 18.6 2.95 ;
      RECT 15.35 1.75 17.5 2 ;
      RECT 16.2 1.05 16.45 2 ;
      RECT 16.35 3.85 16.6 5.3 ;
      RECT 14.65 3.85 14.9 5.3 ;
      RECT 14.65 3.85 16.6 4.1 ;
      RECT 13.75 3.7 14 5.3 ;
      RECT 13.75 3.7 14.3 3.95 ;
      RECT 14.05 2.3 14.3 3.95 ;
      RECT 11.5 2.05 11.8 2.8 ;
      RECT 11.3 2.35 11.8 2.65 ;
      RECT 13.75 2.3 14.3 2.6 ;
      RECT 11.5 2.05 14 2.3 ;
      RECT 13.75 1.05 14 2.6 ;
      RECT 12.35 4.3 12.85 4.6 ;
      RECT 12.45 4.2 12.75 4.6 ;
      RECT 9 2.1 9.3 2.45 ;
      RECT 8.9 2.1 9.4 2.4 ;
      RECT 7.6 4.3 8.15 5.3 ;
      RECT 5.4 4.3 8.15 4.6 ;
      RECT 5.4 2.3 5.7 4.6 ;
      RECT 4.4 3.1 5.7 3.4 ;
      RECT 5.4 2.3 6.55 2.6 ;
      RECT 6.25 1.5 6.55 2.6 ;
      RECT 6.25 1.5 8.15 1.75 ;
      RECT 7.6 1.05 8.15 1.75 ;
      RECT 2.15 1.75 2.4 5.3 ;
      RECT 3.85 2 5.15 2.3 ;
      RECT 3.15 1.7 4.1 2 ;
      RECT 2.15 1.75 4.1 2 ;
      RECT 3.15 1.05 3.4 2 ;
      RECT 4.7 3.85 4.95 5.3 ;
      RECT 3 3.85 3.25 5.3 ;
      RECT 3 3.85 4.95 4.1 ;
      RECT 1.4 1.05 1.65 5.3 ;
      RECT 1.4 2 1.7 2.65 ;
      RECT 1.4 2.3 1.8 2.6 ;
      RECT 16.5 2.25 17 2.55 ;
      RECT 14.6 2.15 15.1 2.45 ;
      RECT 12.35 2.55 12.85 2.85 ;
      RECT 10.7 1.05 11.25 1.95 ;
      RECT 10.7 3.65 11.25 5.3 ;
      RECT 7 2.25 7.5 2.55 ;
      RECT 2.65 2.3 3.15 2.6 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dffsr_1
