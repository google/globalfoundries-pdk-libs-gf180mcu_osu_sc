# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_clkbuf_8
  CLASS CORE ;
  ORIGIN 0.85 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_clkbuf_8 -0.85 -0.15 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.2 4 0.7 4.3 ;
      LAYER MET2 ;
        RECT 0.2 4 0.7 4.3 ;
        RECT 0.25 3.95 0.65 4.35 ;
      LAYER VIA12 ;
        RECT 0.32 4.02 0.58 4.28 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -0.85 7.35 8.15 7.95 ;
        RECT 7.35 5.3 7.6 7.95 ;
        RECT 5.65 5.3 5.9 7.95 ;
        RECT 3.95 5.3 4.2 7.95 ;
        RECT 2.25 5.3 2.5 7.95 ;
        RECT 0.55 5.3 0.8 7.95 ;
      LAYER MET2 ;
        RECT 5.6 7.4 6.1 7.7 ;
        RECT 5.65 7.35 6.05 7.75 ;
        RECT 4.4 7.4 4.9 7.7 ;
        RECT 4.45 7.35 4.85 7.75 ;
        RECT 3.2 7.4 3.7 7.7 ;
        RECT 3.25 7.35 3.65 7.75 ;
        RECT 2 7.4 2.5 7.7 ;
        RECT 2.05 7.35 2.45 7.75 ;
        RECT 0.8 7.4 1.3 7.7 ;
        RECT 0.85 7.35 1.25 7.75 ;
        RECT -0.4 7.4 0.1 7.7 ;
        RECT -0.35 7.35 0.05 7.75 ;
      LAYER VIA12 ;
        RECT -0.28 7.42 -0.02 7.68 ;
        RECT 0.92 7.42 1.18 7.68 ;
        RECT 2.12 7.42 2.38 7.68 ;
        RECT 3.32 7.42 3.58 7.68 ;
        RECT 4.52 7.42 4.78 7.68 ;
        RECT 5.72 7.42 5.98 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -0.85 -0.15 8.15 0.45 ;
        RECT 7.35 -0.15 7.6 1.65 ;
        RECT 5.65 -0.15 5.9 1.65 ;
        RECT 3.95 -0.15 4.2 1.65 ;
        RECT 2.25 -0.15 2.5 1.65 ;
        RECT 0.55 -0.15 0.8 1.65 ;
      LAYER MET2 ;
        RECT 5.6 0.1 6.1 0.4 ;
        RECT 5.65 0.05 6.05 0.45 ;
        RECT 4.4 0.1 4.9 0.4 ;
        RECT 4.45 0.05 4.85 0.45 ;
        RECT 3.2 0.1 3.7 0.4 ;
        RECT 3.25 0.05 3.65 0.45 ;
        RECT 2 0.1 2.5 0.4 ;
        RECT 2.05 0.05 2.45 0.45 ;
        RECT 0.8 0.1 1.3 0.4 ;
        RECT 0.85 0.05 1.25 0.45 ;
        RECT -0.4 0.1 0.1 0.4 ;
        RECT -0.35 0.05 0.05 0.45 ;
      LAYER VIA12 ;
        RECT -0.28 0.12 -0.02 0.38 ;
        RECT 0.92 0.12 1.18 0.38 ;
        RECT 2.12 0.12 2.38 0.38 ;
        RECT 3.32 0.12 3.58 0.38 ;
        RECT 4.52 0.12 4.78 0.38 ;
        RECT 5.72 0.12 5.98 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 4.7 6.9 5 ;
        RECT 6.5 0.8 6.75 7 ;
        RECT 1.4 1.9 6.75 2.15 ;
        RECT 4.8 0.8 5.05 7 ;
        RECT 3.1 0.8 3.35 7 ;
        RECT 1.4 0.8 1.65 7 ;
      LAYER MET2 ;
        RECT 6.4 4.65 6.9 5.05 ;
        RECT 6.35 4.7 6.9 5 ;
      LAYER VIA12 ;
        RECT 6.52 4.72 6.78 4.98 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT -0.3 0.8 -0.05 7 ;
      RECT -0.3 2.75 1.15 3.05 ;
  END
END gf180mcu_osu_sc_12T_clkbuf_8
