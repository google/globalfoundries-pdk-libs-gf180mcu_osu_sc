# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffrn_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffrn_1 0 0 ;
  SIZE 17.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 17.6 8.1 ;
        RECT 15.95 5.45 16.2 8.1 ;
        RECT 12.95 5.45 13.2 8.1 ;
        RECT 10.75 6.2 11 8.1 ;
        RECT 7.95 5.45 8.2 8.1 ;
        RECT 4.9 5.45 5.15 8.1 ;
        RECT 3.55 5.45 3.8 8.1 ;
        RECT 0.55 5.45 0.8 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 17.6 0.6 ;
        RECT 15.95 0 16.2 1.8 ;
        RECT 14.2 0 14.45 1.8 ;
        RECT 12.5 0 12.75 1.8 ;
        RECT 10.75 0 11 1.8 ;
        RECT 7.95 0 8.2 1.4 ;
        RECT 4.9 0 5.15 1.8 ;
        RECT 4 0 4.25 1.8 ;
        RECT 2.3 0 2.55 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 11.15 4.15 11.65 4.45 ;
        RECT 9 4.15 10.05 4.45 ;
        RECT 8.9 2.15 9.4 2.45 ;
        RECT 9 2.15 9.3 4.45 ;
        RECT 6.1 4.15 7.25 4.45 ;
        RECT 6.75 2.2 7.25 2.5 ;
        RECT 6.85 2.2 7.15 4.45 ;
      LAYER MET2 ;
        RECT 6.75 4.15 11.65 4.45 ;
        RECT 11.2 4.1 11.6 4.5 ;
        RECT 9.55 4.1 10.05 4.5 ;
        RECT 6.75 4.1 7.2 4.5 ;
      LAYER VIA12 ;
        RECT 6.87 4.17 7.13 4.43 ;
        RECT 9.67 4.17 9.93 4.43 ;
        RECT 11.27 4.17 11.53 4.43 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.4 3.5 5.9 3.8 ;
      LAYER MET2 ;
        RECT 5.4 3.45 5.9 3.85 ;
      LAYER VIA12 ;
        RECT 5.52 3.52 5.78 3.78 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 16.8 4.8 17.3 5.15 ;
        RECT 16.8 4.75 17.25 5.15 ;
        RECT 16.8 0.95 17.05 7.15 ;
      LAYER MET2 ;
        RECT 16.8 4.8 17.3 5.1 ;
        RECT 16.85 4.75 17.25 5.15 ;
      LAYER VIA12 ;
        RECT 16.92 4.82 17.18 5.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 15.1 4.15 16.55 4.45 ;
        RECT 16.2 2.05 16.45 4.45 ;
        RECT 15.1 2.05 16.45 2.3 ;
        RECT 15.1 4.15 15.35 7.15 ;
        RECT 15.1 0.95 15.35 2.3 ;
      LAYER MET2 ;
        RECT 16.05 4.15 16.55 4.45 ;
        RECT 16.1 4.1 16.5 4.5 ;
      LAYER VIA12 ;
        RECT 16.17 4.17 16.43 4.43 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.55 4.8 1.05 5.1 ;
      LAYER MET2 ;
        RECT 0.55 4.75 1.05 5.15 ;
      LAYER VIA12 ;
        RECT 0.67 4.82 0.93 5.08 ;
    END
  END RN
  OBS
    LAYER MET2 ;
      RECT 15.35 2.8 15.75 3.2 ;
      RECT 15 2.85 15.8 3.15 ;
      RECT 2.65 3.45 3.15 3.85 ;
      RECT 2.75 0.9 3.05 3.85 ;
      RECT 1.3 2.15 1.8 2.55 ;
      RECT 13.75 2.1 14.35 2.5 ;
      RECT 1.3 2.2 3.05 2.5 ;
      RECT 13.75 0.9 14.05 2.5 ;
      RECT 2.75 0.9 14.05 1.2 ;
      RECT 12.4 2.1 12.9 2.5 ;
      RECT 12.4 1.55 12.8 2.5 ;
      RECT 9.3 1.5 9.7 1.9 ;
      RECT 9.25 1.55 12.8 1.85 ;
      RECT 12.45 4.75 12.85 5.15 ;
      RECT 10.25 4.75 10.65 5.15 ;
      RECT 10.2 4.8 12.9 5.1 ;
      RECT 11.55 2.8 11.95 3.2 ;
      RECT 9.6 2.8 10 3.2 ;
      RECT 9.55 2.85 12.05 3.15 ;
      RECT 10.3 3.45 10.7 3.85 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 7.6 2.15 8 2.55 ;
      RECT 3.85 2.15 4.35 2.55 ;
      RECT 3.85 2.2 8.05 2.5 ;
      RECT 14.25 4.75 14.75 5.15 ;
    LAYER VIA12 ;
      RECT 15.42 2.87 15.68 3.13 ;
      RECT 14.37 4.82 14.63 5.08 ;
      RECT 13.97 2.17 14.23 2.43 ;
      RECT 12.52 2.17 12.78 2.43 ;
      RECT 12.52 4.82 12.78 5.08 ;
      RECT 11.62 2.87 11.88 3.13 ;
      RECT 10.37 3.52 10.63 3.78 ;
      RECT 10.32 4.82 10.58 5.08 ;
      RECT 9.67 2.87 9.93 3.13 ;
      RECT 9.37 1.57 9.63 1.83 ;
      RECT 7.67 2.22 7.93 2.48 ;
      RECT 3.97 2.22 4.23 2.48 ;
      RECT 2.77 3.52 3.03 3.78 ;
      RECT 1.42 2.22 1.68 2.48 ;
    LAYER MET1 ;
      RECT 14.35 2.85 14.6 7.15 ;
      RECT 12.5 4.7 12.8 5.2 ;
      RECT 12.5 4.8 14.75 5.1 ;
      RECT 13.35 2.85 15.8 3.15 ;
      RECT 13.35 0.95 13.6 3.15 ;
      RECT 11.6 4.75 11.85 7.15 ;
      RECT 11.6 4.75 12.15 5 ;
      RECT 11.9 3.55 12.15 5 ;
      RECT 11.6 2.75 11.9 3.8 ;
      RECT 11.6 0.95 11.85 3.8 ;
      RECT 10.2 4.8 10.7 5.1 ;
      RECT 10.3 3.5 10.6 5.1 ;
      RECT 10.25 3.5 10.75 3.8 ;
      RECT 9.35 5.95 9.6 7.15 ;
      RECT 8.45 5.95 9.6 6.2 ;
      RECT 8.45 3.45 8.7 6.2 ;
      RECT 8.4 1.6 8.65 3.7 ;
      RECT 8.4 1.6 9.75 1.85 ;
      RECT 9.35 1.55 9.75 1.85 ;
      RECT 9.35 0.95 9.6 1.85 ;
      RECT 7.55 4.8 8.05 5.1 ;
      RECT 7.65 2.2 7.95 5.1 ;
      RECT 7.55 2.2 8.05 2.5 ;
      RECT 6.55 4.95 6.8 7.15 ;
      RECT 4.9 4.95 6.8 5.2 ;
      RECT 4.9 2.25 5.15 5.2 ;
      RECT 3.85 4.15 5.15 4.45 ;
      RECT 4.9 2.25 5.9 2.5 ;
      RECT 5.5 1.55 5.9 2.5 ;
      RECT 5.5 1.55 6.8 1.8 ;
      RECT 6.55 0.95 6.8 1.8 ;
      RECT 2.15 2.5 2.4 7.15 ;
      RECT 2.15 2.5 3.4 2.75 ;
      RECT 3.15 0.95 3.4 2.75 ;
      RECT 3.95 2.15 4.2 2.55 ;
      RECT 3 2.2 4.35 2.5 ;
      RECT 1.4 0.95 1.65 7.15 ;
      RECT 1.3 2.2 1.8 2.5 ;
      RECT 1.4 2.15 1.7 2.5 ;
      RECT 13.85 2.15 14.35 2.45 ;
      RECT 12.4 2.15 12.9 2.45 ;
      RECT 9.55 2.85 10.05 3.15 ;
      RECT 2.65 3.5 3.15 3.8 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffrn_1
