# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__aoi31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__aoi31_1 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 2.3 6.2 2.55 8.1 ;
        RECT 0.6 5.45 0.85 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.85 0 4.1 1.8 ;
        RECT 1.05 0 1.3 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.1 4.8 1.6 5.1 ;
      LAYER MET2 ;
        RECT 1.1 4.75 1.6 5.15 ;
      LAYER VIA12 ;
        RECT 1.22 4.82 1.48 5.08 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.5 2.4 3.8 ;
      LAYER MET2 ;
        RECT 1.9 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.02 3.52 2.28 3.78 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 4.8 3 5.1 ;
      LAYER MET2 ;
        RECT 2.5 4.75 3 5.15 ;
      LAYER VIA12 ;
        RECT 2.62 4.82 2.88 5.08 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.25 3.5 3.75 3.8 ;
      LAYER MET2 ;
        RECT 3.25 3.45 3.75 3.85 ;
      LAYER VIA12 ;
        RECT 3.37 3.52 3.63 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.9 4.8 4.4 5.1 ;
        RECT 4 2.55 4.25 7.15 ;
        RECT 3 2.55 4.25 2.8 ;
        RECT 3 0.95 3.25 2.8 ;
      LAYER MET2 ;
        RECT 3.9 4.75 4.4 5.15 ;
      LAYER VIA12 ;
        RECT 4.02 4.82 4.28 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.15 5.7 3.4 7.15 ;
      RECT 1.45 5.7 1.7 7.15 ;
      RECT 1.45 5.7 3.4 5.95 ;
  END
END gf180mcu_osu_sc_gp12t3v3__aoi31_1
