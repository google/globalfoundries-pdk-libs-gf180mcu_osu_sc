# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_1 0 0 ;
  SIZE 3.85 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 3.85 6.35 ;
        RECT 1.4 3.6 1.75 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 3.85 0.7 ;
        RECT 1.4 0 1.75 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.6 2.3 2.1 2.6 ;
      LAYER Metal2 ;
        RECT 1.6 2.3 2.1 2.6 ;
        RECT 1.65 2.25 2.05 2.65 ;
      LAYER Via1 ;
        RECT 1.72 2.32 1.98 2.58 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.5 2 2.8 2.5 ;
        RECT 0.8 2.3 1.3 2.6 ;
      LAYER Metal2 ;
        RECT 2.4 2.05 2.9 2.45 ;
        RECT 2.4 1.65 2.8 2.45 ;
        RECT 0.9 1.65 2.8 1.95 ;
        RECT 0.8 2.3 1.3 2.6 ;
        RECT 0.85 2.25 1.25 2.65 ;
        RECT 0.9 1.65 1.2 2.65 ;
      LAYER Via1 ;
        RECT 0.92 2.32 1.18 2.58 ;
        RECT 2.52 2.12 2.78 2.38 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.15 1.35 3.4 4.15 ;
        RECT 2.9 3.85 3.2 4.65 ;
        RECT 2.9 3.85 3.15 5.3 ;
        RECT 2.9 1.05 3.15 1.6 ;
      LAYER Metal2 ;
        RECT 2.8 4.2 3.3 4.6 ;
      LAYER Via1 ;
        RECT 2.92 4.27 3.18 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 0.4 3.55 0.9 3.95 ;
      RECT 0.4 3.6 2 3.9 ;
      RECT 1.7 3.1 2 3.9 ;
      RECT 2.4 3.05 2.9 3.45 ;
      RECT 1.7 3.1 2.9 3.4 ;
    LAYER Via1 ;
      RECT 2.52 3.12 2.78 3.38 ;
      RECT 0.52 3.62 0.78 3.88 ;
    LAYER Metal1 ;
      RECT 0.55 3.05 0.8 5.3 ;
      RECT 0.4 3.6 0.9 3.9 ;
      RECT 0.3 1.65 0.55 3.3 ;
      RECT 0.55 1.05 0.8 1.9 ;
      RECT 2.5 3 2.8 3.5 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_1
