* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__nfet_01v8__toxe_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__vth0_slope_spectre = 0.0
.param sky130_fd_pr__nfet_01v8__voff_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__nfet_01v8__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__nfet_01v8__voff_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__nfet_01v8 d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__nfet_01v8.0 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.536077+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.54086565
+ k2 = -0.030899431
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1814466+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.30474
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.03243309
+ ua = -7.5866357e-10
+ ub = 1.674192e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.297743
+ ags = 0.430444
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -0.0020233
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.1 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.536077+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.54086565
+ k2 = -0.030899431
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.1814466+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.30474
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.03243309
+ ua = -7.5866357e-10
+ ub = 1.674192e-18
+ uc = 4.9242e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.297743
+ ags = 0.430444
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 2.1073424e-24
+ keta = -0.0087946
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.026316
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0030734587
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 754674160.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31303
+ kt2 = -0.045313337
+ at = 140000.0
+ ute = -1.8134
+ ua1 = 3.7602e-10
+ ub1 = -6.3962e-19
+ uc1 = 1.5829713e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -0.0020233
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.2 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.367912299e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(1))} lvth0 = -5.696795150e-09 wvth0 = -7.139176946e-08 pvth0 = 5.694304625e-13
+ k1 = 5.415457968e-01 lk1 = -5.424943089e-09 wk1 = -6.798494173e-08 pk1 = 5.422571412e-13
+ k2 = -3.140779186e-02 lk2 = 4.054755328e-09 wk2 = 5.081386112e-08 pk2 = -4.052982670e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.807326273e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.694743212e-09 wvoff = -7.136605475e-08 pvoff = 5.692253584e-13
+ nfactor = 2.305958637e+00 lnfactor = -9.720015876e-09 wnfactor = -1.218104415e-07 pnfactor = 9.715766479e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.241770275e-02 lu0 = 1.227307679e-10 wu0 = 1.538051914e-09 pu0 = -1.226771124e-14
+ ua = -7.582789781e-10 lua = -3.067557542e-18 wua = -3.844237946e-17 pua = 3.066216468e-22
+ ub = 1.672091096e-18 lub = 1.675709387e-26 wub = 2.099985257e-25 pub = -1.674976801e-30
+ uc = 4.877008480e-11 luc = 3.764059839e-18 wuc = 4.717088911e-17 puc = -3.762414268e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.289305555e+00 la0 = 6.729821120e-08 wa0 = 8.433756617e-07 pa0 = -6.726878977e-12
+ ags = 4.320303102e-01 lags = -1.265262591e-08 wags = -1.585616699e-07 pags = 1.264709444e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.950656262e-24 lb1 = 1.249749944e-30 wb1 = 1.566176377e-29 pb1 = -1.249203578e-34
+ keta = -8.288058846e-03 lketa = -4.040241132e-09 wketa = -5.063197041e-08 pketa = 4.038474820e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.800573404e-02 lpclm = -3.325229885e-07 wpclm = -4.167150812e-06 ppclm = 3.323776161e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.074732157e-03 lpdiblc2 = -1.015726833e-11 wpdiblc2 = -1.272900534e-10 ppdiblc2 = 1.015282777e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.580442487e+08 lpscbe1 = -2.688028581e+01 wpscbe1 = -3.368615365e+02 ppscbe1 = 2.686853428e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.131868837e-01 lkt1 = 1.251326022e-09 wkt1 = 1.568151505e-08 pkt1 = -1.250778967e-13
+ kt2 = -4.539671736e-02 lkt2 = 6.650530936e-10 wkt2 = 8.334390809e-09 pkt2 = -6.647623457e-14
+ at = 140000.0
+ ute = -1.816359229e+00 lute = 2.360321122e-08 wute = 2.957935066e-07 pute = -2.359289237e-12
+ ua1 = 3.613755352e-10 lua1 = 1.168062433e-16 wua1 = 1.463806258e-15 pua1 = -1.167551779e-20
+ ub1 = -6.204482125e-19 lub1 = -1.529167842e-25 wub1 = -1.916340595e-24 pub1 = 1.528499321e-29
+ uc1 = 1.690988400e-11 luc1 = -8.615590785e-18 wuc1 = -1.079698769e-16 puc1 = 8.611824221e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.065673479e-03 ltvoff = 3.379766350e-10 wtvoff = 4.235495463e-09 ptvoff = -3.378288784e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.3 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.257881703e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.805286631e-08 wvth0 = 7.970998398e-08 pvth0 = -3.137065901e-14
+ k1 = 5.304574419e-01 lk1 = 3.866386370e-08 wk1 = 1.369158390e-07 pk1 = -2.724562297e-13
+ k2 = -2.326625831e-02 lk2 = -2.831708931e-08 wk2 = -8.771961924e-08 pk2 = 1.455296915e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.378281302e-01 ldsub = 8.815836977e-08 wdsub = 2.216217672e-06 pdsub = -8.811982869e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.918053716e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.833199408e-08 wvoff = 8.704284409e-08 pvoff = -6.062996693e-14
+ nfactor = 2.285160074e+00 lnfactor = 7.297789931e-08 wnfactor = 3.384011255e-07 pnfactor = -8.582871314e-13
+ eta0 = 7.412445450e-02 leta0 = 2.336196799e-08 weta0 = 5.872976830e-07 peta0 = -2.335175460e-12
+ etab = -6.486356790e-02 letab = -2.042315258e-08 wetab = -5.134186554e-07 petab = 2.041422399e-12
+ u0 = 3.254619738e-02 lu0 = -3.881813322e-10 wu0 = 9.133334821e-09 pu0 = -4.246758904e-14
+ ua = -7.772766349e-10 lua = 7.246970951e-17 wua = 1.349633081e-15 pua = -5.212555164e-21
+ ub = 1.715448650e-18 lub = -1.556384353e-25 wub = -1.333196930e-24 pub = 4.460978208e-30
+ uc = 5.877915793e-11 luc = -3.603337616e-17 wuc = -3.264462550e-16 puc = 1.109311150e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.424425234e+00 la0 = -4.699560085e-07 wa0 = -1.455090090e-06 pa0 = 2.412133444e-12
+ ags = 4.202144348e-01 lags = 3.432890182e-08 wags = -1.084612175e-06 pags = 4.946812196e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 4.502912266e-24 lb1 = -8.898367034e-30 wb1 = -3.132352754e-29 pb1 = 6.189955043e-35
+ keta = -1.640202815e-02 lketa = 2.822200432e-08 wketa = 8.756343093e-08 pketa = -1.456362283e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.131369147e-01 lpclm = 2.375792818e-06 wpclm = 8.540188246e-06 ppclm = -1.728834668e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.181248537e-03 lpdiblc2 = -4.336808822e-10 wpdiblc2 = -1.246582526e-08 ppdiblc2 = 5.007497679e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.031489705e+08 lpscbe1 = 1.913908060e+02 wpscbe1 = 6.737230730e+02 ppscbe1 = -1.331368419e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.112847401e-01 lkt1 = -6.311855597e-09 wkt1 = 3.394151730e-08 pkt1 = -1.976821490e-13
+ kt2 = -4.403955904e-02 lkt2 = -4.731192969e-09 wkt2 = -1.656662876e-08 pkt2 = 3.253360577e-14
+ at = 1.381479098e+05 lat = 7.364162488e-03 wat = 1.851280495e-01 pat = -7.360943023e-7
+ ute = -1.757935204e+00 lute = -2.086986568e-07 wute = -1.613263360e-06 pute = 5.231380497e-12
+ ua1 = 6.225548039e-10 lua1 = -9.216780498e-16 wua1 = -5.190223011e-15 pua1 = 1.478180753e-20
+ ub1 = -9.463016587e-19 lub1 = 1.142720834e-24 wub1 = 5.188563162e-24 pub1 = -1.296507040e-29
+ uc1 = -2.357426518e-13 luc1 = 5.955775258e-17 wuc1 = 1.710346184e-16 puc1 = -2.481773957e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.421023671e-03 ltvoff = -2.225238676e-09 wtvoff = -3.915924870e-09 ptvoff = -1.371732000e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.4 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.461881904e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.260347812e-09 wvth0 = -5.049695639e-08 pvth0 = 2.259359633e-13
+ k1 = 5.524870904e-01 lk1 = -4.869717742e-09 wk1 = -2.472758915e-07 pk1 = 4.867588799e-13
+ k2 = -3.838702190e-02 lk2 = 1.563595979e-09 wk2 = 6.501325548e-08 pk2 = -1.562912406e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 5.824396194e-01 wdsub = -2.242980920e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.731593458e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.484911228e-09 wvoff = 1.314710811e-07 pvoff = -1.484262055e-13
+ nfactor = 2.306233618e+00 lnfactor = 3.133371024e-08 wnfactor = 1.488986938e-06 pnfactor = -3.132001177e-12
+ eta0 = 8.609480828e-02 leta0 = -2.930790459e-10 weta0 = -6.092143748e-07 peta0 = 2.929509176e-14
+ etab = -7.518471959e-02 letab = -2.715316148e-11 wetab = 5.182452938e-07 petab = 2.714129066e-15
+ u0 = 3.203839579e-02 lu0 = 6.153036758e-10 wu0 = 1.876621368e-08 pu0 = -6.150346773e-14
+ ua = -7.784147269e-10 lua = 7.471873419e-17 wua = 2.491281076e-15 pua = -7.468606865e-21
+ ub = 1.671533075e-18 lub = -6.885528766e-26 wub = -2.558588474e-24 pub = 6.882518551e-30
+ uc = 3.956352106e-11 luc = 1.939335609e-18 wuc = 3.330022481e-16 puc = -1.938487771e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.148217881e+04 lvsat = -2.928986896e-03 wvsat = -1.481530827e-01 pvsat = 2.927706402e-7
+ a0 = 1.176203689e+00 la0 = 2.056352243e-08 wa0 = 8.056787490e-07 pa0 = -2.055453247e-12
+ ags = 4.608595850e-01 lags = -4.599144281e-08 wags = -9.076615155e-07 pags = 4.597133627e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.862460185e-03 lketa = 9.370520639e-09 wketa = 4.878426501e-07 pketa = -9.366424034e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.768770306e-01 lpclm = 2.416342047e-08 wpclm = 1.013853514e-06 ppclm = -2.415285670e-12
+ pdiblc1 = 4.131572185e-01 lpdiblc1 = -4.576181312e-08 wpdiblc1 = -2.314709462e-06 ppdiblc1 = 4.574180697e-12
+ pdiblc2 = 2.903299932e-03 lpdiblc2 = 1.155833635e-10 wpdiblc2 = 1.872041904e-08 ppdiblc2 = -1.155328327e-14
+ pdiblcb = -2.318864550e-02 lpdiblcb = -3.579482830e-09 wpdiblcb = -1.810562609e-07 ppdiblcb = 3.577917952e-13
+ drout = 5.380958797e-01 ldrout = 4.328552063e-08 wdrout = 2.189454424e-06 pdrout = -4.326659707e-12
+ pscbe1 = 7.606510411e+08 lpscbe1 = 7.775889417e+01 wpscbe1 = 3.933175629e+03 ppscbe1 = -7.772489954e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.205658464e-07 lalpha0 = -3.765840295e-13 walpha0 = -1.904825348e-11 palpha0 = 3.764193945e-17
+ alpha1 = 8.524824670e-01 lalpha1 = -4.905692338e-09 walpha1 = -2.481381680e-07 palpha1 = 4.903547668e-13
+ beta0 = 1.406239407e+01 lbeta0 = -3.999582106e-07 wbeta0 = -2.023055887e-05 pbeta0 = 3.997833569e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.107339048e-01 lkt1 = -7.400381177e-09 wkt1 = -4.404168957e-07 pkt1 = 7.397145879e-13
+ kt2 = -4.496893626e-02 lkt2 = -2.894617183e-09 wkt2 = -1.465179912e-07 pkt2 = 2.893351714e-13
+ at = 1.381088459e+05 lat = 7.441358137e-03 wat = 1.890327353e-01 pat = -7.438104924e-7
+ ute = -1.803083395e+00 lute = -1.194796923e-07 wute = -5.009469552e-06 pute = 1.194274582e-11
+ ua1 = 2.816514627e-10 lua1 = -2.480066846e-16 wua1 = -1.025466117e-14 pua1 = 2.478982610e-20
+ ub1 = -4.339323422e-19 lub1 = 1.302093822e-25 wub1 = 5.213953787e-24 pub1 = -1.301524572e-29
+ uc1 = 3.132149136e-11 luc1 = -2.803633615e-18 wuc1 = -9.636508894e-17 puc1 = 2.802407923e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.537784454e-03 ltvoff = -1.836748925e-11 wtvoff = -5.539131945e-09 ptvoff = 1.835945936e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.5 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.364286978e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.266244272e-09 wvth0 = 1.123312552e-07 pvth0 = 6.699348414e-14
+ k1 = 5.406566785e-01 lk1 = 6.678373256e-09 wk1 = 9.474366135e-07 pk1 = -6.794430059e-13
+ k2 = -3.211294494e-02 lk2 = -4.560756409e-09 wk2 = -3.829160891e-07 pk2 = 2.809487180e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.991414420e-01 ldsub = -3.091440504e-07 wdsub = -5.343647045e-06 pdsub = 3.026671828e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.807804359e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 8.924131638e-09 wvoff = 1.756981189e-07 pvoff = -1.915978092e-13
+ nfactor = 2.359007702e+00 lnfactor = -2.018097312e-08 wnfactor = -2.564883450e-06 pnfactor = 8.251276484e-13
+ eta0 = 2.018846564e-01 leta0 = -1.133197182e-07 weta0 = -4.615884383e-06 peta0 = 3.940349927e-12
+ etab = -1.463451305e-01 letab = 6.943508571e-08 wetab = 1.015844159e-06 petab = -4.830100369e-13
+ u0 = 3.419554615e-02 lu0 = -1.490368454e-09 wu0 = -3.953752008e-08 pu0 = -4.591094276e-15
+ ua = -5.371888159e-10 lua = -1.607505616e-16 wua = -5.221570888e-15 pua = 6.018559916e-23
+ ub = 1.475966341e-18 lub = 1.220444419e-25 wub = 5.223075908e-24 pub = -7.134441927e-31
+ uc = 1.095109860e-11 luc = 2.986895122e-17 wuc = 2.023582373e-16 puc = -6.632245490e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.966833487e+04 lvsat = -1.158428535e-03 wvsat = 3.315201299e-02 pvsat = 1.157922093e-7
+ a0 = 1.264240561e+00 la0 = -6.537243798e-08 wa0 = -5.009235444e-06 pa0 = 3.620693833e-12
+ ags = 2.401739658e-01 lags = 1.694277348e-07 wags = 3.090076394e-06 pags = 6.947977349e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 3.561401696e-03 lketa = -8.045862015e-10 wketa = -7.306170793e-07 pketa = 2.527400029e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.404786183e-01 lpclm = -3.792037900e-08 wpclm = -2.690702931e-06 ppclm = 1.200865240e-12
+ pdiblc1 = 3.871350928e-01 lpdiblc1 = -2.036067943e-08 wpdiblc1 = 2.863654728e-07 ppdiblc1 = 2.035177815e-12
+ pdiblc2 = 1.217587306e-03 lpdiblc2 = 1.761068143e-09 wpdiblc2 = 2.331725074e-08 ppdiblc2 = -1.604041618e-14
+ pdiblcb = -2.862270899e-02 lpdiblcb = 1.724902169e-09 wpdiblcb = 3.621125218e-07 ppdiblcb = -1.724148077e-13
+ drout = 5.994456506e-01 ldrout = -1.660019935e-08 wdrout = -3.942840578e-06 pdrout = 1.659294207e-12
+ pscbe1 = 8.616614397e+08 lpscbe1 = -2.084099226e+01 wpscbe1 = -6.163448258e+03 ppscbe1 = 2.083188100e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.410386908e-08 lalpha0 = -2.336172208e-13 walpha0 = -4.408458775e-12 palpha0 = 2.335150880e-17
+ alpha1 = 8.450350661e-01 lalpha1 = 2.363983782e-09 walpha1 = 4.962763360e-07 palpha1 = -2.362950295e-13
+ beta0 = 1.380708182e+01 lbeta0 = -1.507387305e-07 wbeta0 = 5.289504551e-06 pbeta0 = 1.506728306e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.095566483e-01 lkt1 = -8.549543620e-09 wkt1 = 2.833493486e-07 pkt1 = 3.322030121e-14
+ kt2 = -4.861045418e-02 lkt2 = 6.599995580e-10 wkt2 = 2.187908274e-07 pkt2 = -6.725591757e-14
+ at = 1.706731833e+05 lat = -2.434586389e-02 wat = -6.806270065e-01 pat = 1.050956893e-7
+ ute = -2.105517726e+00 lute = 1.757373462e-07 wute = 1.205657763e-05 pute = -4.716037219e-12
+ ua1 = -3.629341746e-10 lua1 = 3.811965610e-16 wua1 = 2.502228661e-14 pua1 = -9.645272601e-21
+ ub1 = -9.356348756e-20 lub1 = -2.020369101e-25 wub1 = -1.133769218e-23 pub1 = 3.141411760e-30
+ uc1 = 1.727110250e-11 luc1 = 1.091145677e-17 wuc1 = 7.294628321e-16 puc1 = -5.258795712e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.890636836e-03 ltvoff = -6.500715761e-10 wtvoff = -1.153418012e-08 ptvoff = 7.687928284e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.6 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.487389318e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.404898722e-09 wvth0 = 5.479671596e-07 pvth0 = -1.404284528e-13
+ k1 = 5.733572999e-01 lk1 = -8.891569812e-09 wk1 = -2.346183834e-06 pk1 = 8.887682595e-13
+ k2 = -4.702258562e-02 lk2 = 2.538260265e-09 wk2 = 7.400063047e-07 pk2 = -2.537150589e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.608544335e-01 ldsub = -5.232627283e-09 wdsub = -8.540599614e-08 pdsub = 5.230339683e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.633755034e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 6.370166662e-10 wvoff = -9.297299967e-08 pvoff = -6.367381753e-14
+ nfactor = 2.331268357e+00 lnfactor = -6.973272136e-09 wnfactor = -2.295831557e-06 pnfactor = 6.970223560e-13
+ eta0 = -3.611397891e-02 weta0 = 3.659797201e-6
+ etab = -5.538291750e-04 letab = 1.859865862e-11 wetab = 5.311487409e-09 petab = -1.859052765e-15
+ u0 = 3.066008519e-02 lu0 = 1.929917864e-10 wu0 = -8.664729230e-09 pu0 = -1.929074142e-14
+ ua = -9.104153604e-10 lua = 1.695603236e-17 wua = -1.535549350e-15 pua = -1.694861952e-21
+ ub = 1.754640735e-18 lub = -1.064246927e-26 wub = 1.490474610e-24 pub = 1.063781659e-30
+ uc = 7.380749713e-11 luc = -5.924295007e-20 wuc = 5.062814353e-17 puc = 5.921705023e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.890265507e+04 lvsat = -7.938608141e-04 wvsat = 1.096865197e-01 pvsat = 7.935137540e-8
+ a0 = 1.126942734e+00 wa0 = 2.595091542e-6
+ ags = 5.127609304e-01 lags = 3.963926782e-08 wags = 1.287087761e-05 pags = -3.962193833e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.079528043e-03 lketa = 3.771231919e-10 wketa = -1.206320433e-07 pketa = -3.769583212e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.524057554e-01 lpclm = 4.014281679e-09 wpclm = 6.741296190e-07 ppclm = -4.012526715e-13
+ pdiblc1 = 2.847083853e-01 lpdiblc1 = 2.840836336e-08 wpdiblc1 = 1.052455833e-05 ppdiblc1 = -2.839594379e-12
+ pdiblc2 = 4.856343117e-03 lpdiblc2 = 2.852550623e-11 wpdiblc2 = -4.383054714e-09 ppdiblc2 = -2.851303545e-15
+ pdiblcb = -3.853174870e-02 lpdiblcb = 6.442952699e-09 wpdiblcb = 1.352583289e-06 ppdiblcb = -6.440135969e-13
+ drout = 5.984950270e-01 ldrout = -1.614757321e-08 wdrout = -3.847819773e-06 pdrout = 1.614051381e-12
+ pscbe1 = 8.340729560e+08 lpscbe1 = -7.705121978e+00 wpscbe1 = -3.405805999e+03 ppscbe1 = 7.701753453e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.438818033e-07 lalpha0 = 1.082416053e-13 walpha0 = 6.735871957e-11 palpha0 = -1.081942843e-17
+ alpha1 = 0.85
+ beta0 = 1.351261868e+01 lbeta0 = -1.053422766e-08 wbeta0 = 3.472294548e-05 pbeta0 = 1.052962231e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.285216740e-01 lkt1 = 4.803878418e-10 wkt1 = 4.539688434e-07 pkt1 = -4.801778259e-14
+ kt2 = -4.748635604e-02 lkt2 = 1.247759616e-10 wkt2 = 1.037317342e-07 pkt2 = -1.247214120e-14
+ at = 1.176801617e+05 lat = 8.860214216e-04 wat = -2.738963741e-01 pat = -8.856340708e-8
+ ute = -1.698659221e+00 lute = -1.798263502e-08 wute = -1.623367921e-06 pute = 1.797477337e-12
+ ua1 = 4.605278602e-10 lua1 = -1.088335838e-17 wua1 = 2.480129244e-15 pua1 = 1.087860040e-21
+ ub1 = -4.886624463e-19 lub1 = -1.391607233e-26 wub1 = -7.661404497e-24 pub1 = 1.390998850e-30
+ uc1 = 4.720982253e-11 luc1 = -3.343445632e-18 wuc1 = -1.076907545e-15 puc1 = 3.341983944e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.259996096e-03 ltvoff = 1.929664333e-12 wtvoff = 5.017415127e-09 ptvoff = -1.928820723e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.7 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.467620854e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.851934849e-09 wvth0 = 7.455653714e-07 pvth0 = -1.851125220e-13
+ k1 = 5.548884107e-01 lk1 = -4.715089080e-09 wk1 = -5.001023353e-07 pk1 = 4.713027737e-13
+ k2 = -4.250827421e-02 lk2 = 1.517411939e-09 wk2 = 2.887725198e-07 pk2 = -1.516748557e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.111893909e-01 ldsub = 5.998426783e-09 wdsub = 4.878927004e-06 pdsub = -5.995804390e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.668102889e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.413745330e-09 wvoff = 2.503553928e-07 pvoff = -1.413127269e-13
+ nfactor = 2.313012670e+00 lnfactor = -2.845004206e-09 wnfactor = -4.710610058e-07 pnfactor = 2.843760427e-13
+ eta0 = -1.126962478e-01 leta0 = 1.731800795e-08 weta0 = 1.131467606e-05 peta0 = -1.731043687e-12
+ etab = -5.054282121e-03 letab = 1.036313086e-09 wetab = 4.551600312e-07 petab = -1.035860031e-13
+ u0 = 3.361630265e-02 lu0 = -4.755154051e-10 wu0 = -3.041572353e-07 pu0 = 4.753075193e-14
+ ua = -6.073824236e-10 lua = -5.157062385e-17 wua = -3.182559504e-14 pua = 5.154807821e-21
+ ub = 1.544202603e-18 lub = 3.694516816e-26 wub = 2.252508788e-23 pub = -3.692901647e-30
+ uc = 7.384766442e-11 luc = -6.832622020e-20 wuc = 4.661317063e-17 puc = 6.829634934e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.743615097e+04 lvsat = -4.622314448e-04 wvsat = 2.562728163e-01 pvsat = 4.620293665e-8
+ a0 = 1.126942734e+00 wa0 = 2.595091542e-6
+ ags = 8.933414399e-01 lags = -4.642368628e-08 wags = -2.517053512e-05 pags = 4.640339077e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.632681265e-03 lketa = 2.589933484e-11 wketa = -2.758794648e-07 pketa = -2.588801217e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.492089963e-01 lpclm = 4.737183991e-09 wpclm = 9.936657716e-07 ppclm = -4.735112989e-13
+ pdiblc1 = 4.531641189e-01 lpdiblc1 = -9.685542409e-09 wpdiblc1 = -6.313650481e-06 ppdiblc1 = 9.681308084e-13
+ pdiblc2 = 6.031854250e-03 lpdiblc2 = -2.372998792e-10 wpdiblc2 = -1.218827769e-07 ppdiblc2 = 2.371961364e-14
+ pdiblcb = 1.309104138e-02 lpdiblcb = -5.230818559e-09 wpdiblcb = -3.807438874e-06 ppdiblcb = 5.228531750e-13
+ drout = 4.798565019e-01 ldrout = 1.068086830e-08 wdrout = 8.010846098e-06 pdrout = -1.067619884e-12
+ pscbe1 = 7.993153719e+08 lpscbe1 = 1.548190656e-01 wpscbe1 = 6.843288191e+01 ppscbe1 = -1.547513818e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.040459718e-07 lalpha0 = 9.923328974e-14 walpha0 = 6.337687796e-11 palpha0 = -9.918990693e-18
+ alpha1 = 9.069090007e-01 lalpha1 = -1.286917378e-08 walpha1 = -5.688412120e-06 palpha1 = 1.286354763e-12
+ beta0 = 1.277748789e+01 lbeta0 = 1.557053069e-07 wbeta0 = 1.082038852e-04 pbeta0 = -1.556372356e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.209694650e-01 lkt1 = -1.227438479e-09 wkt1 = -3.009218830e-07 pkt1 = 1.226901867e-13
+ kt2 = -4.630223396e-02 lkt2 = -1.429966677e-10 wkt2 = -1.462870566e-08 pkt2 = 1.429341524e-14
+ at = 1.232736586e+05 lat = -3.788696079e-04 wat = -8.330015340e-01 pat = 3.787039736e-8
+ ute = -1.937606266e+00 lute = 3.605189395e-08 wute = 2.226089029e-05 pute = -3.603613278e-12
+ ua1 = 7.614258198e-11 lua1 = 7.603999089e-17 wua1 = 4.090185251e-14 pua1 = -7.600674773e-21
+ ub1 = -2.691863256e-19 lub1 = -6.354752435e-26 wub1 = -2.959942151e-23 pub1 = 6.351974265e-30
+ uc1 = 3.935986943e-11 luc1 = -1.568288639e-18 wuc1 = -2.922554192e-16 puc1 = 1.567603014e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.974350596e-03 ltvoff = -6.266506651e-11 wtvoff = -2.353464705e-08 ptvoff = 6.263767059e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.8 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.0e-06 wmax = 0.0001
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.421562290e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.571074836e-09 wvth0 = 1.205949647e-06 pvth0 = -2.569950814e-13
+ k1 = 5.297223808e-01 lk1 = -7.857658419e-10 wk1 = 2.015400442e-06 pk1 = 7.854223208e-14
+ k2 = -3.293978270e-02 lk2 = 2.342594867e-11 wk2 = -6.676583159e-07 pk2 = -2.341570731e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.268343873e-01 ldsub = 3.555679632e-09 wdsub = 3.315111336e-06 pdsub = -3.554125160e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.701734074e-03 lcdscd = 2.651605064e-10 wcdscd = 1.697523848e-07 pcdscd = -2.650445835e-14
+ cit = 0.0
+ voff = {-1.596489650e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.956048609e-10 wvoff = -4.654639189e-07 pvoff = -2.954756283e-14
+ nfactor = 2.237811370e+00 lnfactor = 8.896626028e-09 wnfactor = 7.045781381e-06 pnfactor = -8.892736601e-13
+ eta0 = -1.127808870e-02 leta0 = 1.482982266e-09 weta0 = 1.177293955e-06 peta0 = -1.482333935e-13
+ etab = -2.892433920e-03 letab = 6.987707553e-10 wetab = 2.390697228e-07 petab = -6.984652667e-14
+ u0 = 2.637508936e-02 lu0 = 6.550986726e-10 wu0 = 4.196475220e-07 pu0 = -6.548122766e-14
+ ua = -1.451257292e-09 lua = 8.018862258e-17 wua = 5.252499926e-14 pua = -8.015356571e-21
+ ub = 2.213250091e-18 lub = -6.751723050e-26 wub = -4.435041155e-23 pub = 6.748771332e-30
+ uc = 6.294653549e-11 luc = 1.633732446e-18 wuc = 1.136249488e-15 puc = -1.633018211e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.823516818e+04 lvsat = -5.869867951e-04 wvsat = 1.764060272e-01 pvsat = 5.867301762e-8
+ a0 = 1.126942734e+00 wa0 = 2.595091542e-6
+ ags = 5.960129168e-01 wags = 4.549318575e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.221854762e-02 lketa = -3.032159495e-09 wketa = -2.233609846e-06 pketa = 3.030833895e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.427722098e-01 lpclm = 5.742198078e-09 wpclm = 1.637063011e-06 ppclm = -5.739687704e-13
+ pdiblc1 = 3.948535541e-01 lpdiblc1 = -5.811640668e-10 wpdiblc1 = -4.851432247e-07 ppdiblc1 = 5.809099935e-14
+ pdiblc2 = 4.739215410e-03 lpdiblc2 = -3.547242126e-11 wpdiblc2 = 7.324595465e-09 ppdiblc2 = 3.545691343e-15
+ pdiblcb = 6.744804231e-03 lpdiblcb = -4.239942475e-09 wpdiblcb = -3.173092604e-06 ppdiblcb = 4.238088857e-13
+ drout = 4.915551465e-01 ldrout = 8.854288734e-09 wdrout = 6.841493081e-06 pdrout = -8.850417816e-13
+ pscbe1 = 7.986209646e+08 lpscbe1 = 2.632410390e-01 wpscbe1 = 1.378432507e+02 ppscbe1 = -2.631259553e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.786292971e-08 lalpha0 = -9.917985016e-16 walpha0 = -7.859492192e-13 palpha0 = 9.913649071e-20
+ alpha1 = 7.172123318e-01 lalpha1 = 1.674930532e-08 walpha1 = 1.327296161e-05 palpha1 = -1.674198286e-12
+ beta0 = 1.341620656e+01 lbeta0 = 5.597832913e-08 wbeta0 = 4.435994207e-05 pbeta0 = -5.595385653e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.150847439e-01 lkt1 = -2.146255297e-09 wkt1 = -8.891367274e-07 pkt1 = 2.145316997e-13
+ kt2 = -4.510229766e-02 lkt2 = -3.303499223e-10 wkt2 = -1.345698772e-07 pkt2 = 3.302054999e-14
+ at = 1.198289709e+05 lat = 1.589701562e-04 wat = -4.886833555e-01 pat = -1.589006576e-8
+ ute = -1.132927038e+00 lute = -8.958750189e-08 wute = -5.817185347e-05 pute = 8.954833602e-12
+ ua1 = 1.362272965e-09 lua1 = -1.247712625e-16 wua1 = -8.765495871e-14 pua1 = 1.247167150e-20
+ ub1 = -1.134148121e-18 lub1 = 7.150415049e-26 wub1 = 5.685894360e-23 pub1 = -7.147289030e-30
+ uc1 = 3.786297182e-11 luc1 = -1.334569033e-18 wuc1 = -1.426310994e-16 puc1 = 1.333985586e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.553247297e-03 ltvoff = 2.772154887e-11 wtvoff = 3.432971489e-08 ptvoff = -2.770942956e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.9 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.371883577e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.111092438e-07 wvth0 = -7.730917236e-09 pvth0 = 7.729072330e-13
+ k1 = 5.418171603e-01 lk1 = -9.512831965e-08 wk1 = -6.618973728e-09 pk1 = 6.617394176e-13
+ k2 = -3.129196426e-02 lk2 = 3.924395815e-08 wk2 = 2.730572021e-09 pk2 = -2.729920397e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.956627950e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.421280247e-06 wvoff = 9.889186155e-08 pvoff = -9.886826200e-12
+ nfactor = 2.387955689e+00 lnfactor = -8.319583025e-06 wnfactor = -5.788717984e-07 pnfactor = 5.787336564e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.216410556e-02 lu0 = 2.689202517e-08 wu0 = 1.871131633e-09 pu0 = -1.870685106e-13
+ ua = -7.362717244e-10 lua = -2.238650203e-15 wua = -1.557639926e-16 pua = 1.557268211e-20
+ ub = 1.621184695e-18 lub = 5.299465505e-24 wub = 3.687337596e-25 pub = -3.686457650e-29
+ uc = 4.772038059e-11 luc = 1.521256295e-16 wuc = 1.058481374e-17 puc = -1.058228778e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.309677100e+00 la0 = -1.193125210e-06 wa0 = -8.301696538e-08 pa0 = 8.299715421e-12
+ ags = 4.288704017e-01 lags = 1.573222757e-07 wags = 1.094639339e-08 pags = -1.094378114e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 8.033273090e-25 lb1 = 1.303703901e-28 wb1 = 9.071096705e-30 pb1 = -9.068931979e-34
+ keta = -7.180997052e-03 lketa = -1.613217878e-07 wketa = -1.122467714e-08 pketa = 1.122199848e-12
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.760603957e-02 lpclm = -3.128257252e-06 wpclm = -2.176623391e-07 ppclm = 2.176103961e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.147856669e-03 lpdiblc2 = -7.438021498e-09 wpdiblc2 = -5.175332547e-10 ppdiblc2 = 5.174097506e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.174573788e+08 lpscbe1 = 3.720789982e+03 wpscbe1 = 2.588904254e+02 ppscbe1 = -2.588286437e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.200657108e-01 lkt1 = 7.034031752e-07 wkt1 = 4.894238807e-08 pkt1 = -4.893070846e-12
+ kt2 = -4.543472374e-02 lkt2 = 1.213577724e-08 wkt2 = 8.444003956e-10 pkt2 = -8.441988879e-14
+ at = 140000.0
+ ute = -1.856901360e+00 lute = 4.349097908e-06 wute = 3.026077292e-07 pute = -3.025355149e-11
+ ua1 = 3.036703693e-10 lua1 = 7.233236521e-15 wua1 = 5.032844339e-16 pua1 = -5.031643301e-20
+ ub1 = -5.518932882e-19 lub1 = -8.770577673e-24 wub1 = -6.102517464e-25 pub1 = 6.101061160e-29
+ uc1 = 1.657054426e-11 luc1 = -7.406544670e-17 wuc1 = -5.153431152e-18 puc1 = 5.152201337e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.344103300e-03 ltvoff = -6.790346166e-08 wtvoff = -4.724683779e-09 ptvoff = 4.723556281e-13
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.10 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.316262588e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} wvth0 = 3.096061115e-8
+ k1 = 5.370550621e-01 wk1 = 2.650752369e-8
+ k2 = -2.932742226e-02 wk2 = -1.093533613e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.245138878e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} wvoff = -3.960400011e-7
+ nfactor = 1.971479598e+00 wnfactor = 2.318253334e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.351031311e-02 wu0 = -7.493467739e-9
+ ua = -8.483379519e-10 wua = 6.238002890e-16
+ ub = 1.886474514e-18 wub = -1.476697033e-24
+ uc = 5.533574872e-11 wuc = -4.238983453e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.249949573e+00 wa0 = 3.324645582e-7
+ ags = 4.367459126e-01 wags = -4.383788093e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 7.329634002e-24 wb1 = -3.632773307e-29
+ keta = -1.525672240e-02 wketa = 4.495234571e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.899367781e-02 wpclm = 8.716894561e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 2.775511312e-03 wpdiblc2 = 2.072606052e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 9.037191254e+08 wpscbe1 = -1.036798810e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.848535368e-01 wkt1 = -1.960034236e-7
+ kt2 = -4.482720999e-02 wkt2 = -3.381636551e-9
+ at = 140000.0
+ ute = -1.639186688e+00 wute = -1.211876929e-6
+ ua1 = 6.657642457e-10 wua1 = -2.015542681e-15
+ ub1 = -9.909460496e-19 wub1 = 2.443923075e-24
+ uc1 = 1.286284790e-11 wuc1 = 2.063835029e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.743332343e-03 wtvoff = 1.892131203e-8
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.11 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.179563729e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.090328689e-07 wvth0 = 5.962880766e-08 pvth0 = -2.286614343e-13
+ k1 = 5.247112438e-01 lk1 = 9.845597383e-08 wk1 = 4.912095597e-08 pk1 = -1.803678113e-13
+ k2 = -1.968728600e-02 lk2 = -7.689103782e-08 wk2 = -3.071728278e-08 pk2 = 1.577834969e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.255062917e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.915548373e-09 wvoff = -4.555360193e-07 pvoff = 4.745483321e-13
+ nfactor = 1.923631785e+00 lnfactor = 3.816406629e-07 wnfactor = 2.537762955e-06 pnfactor = -1.750838597e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.464606866e-02 lu0 = -9.058940723e-09 wu0 = -1.396308973e-08 pu0 = 5.160258488e-14
+ ua = -8.875308152e-10 lua = 3.126076079e-16 wua = 8.606698490e-16 pua = -1.889303825e-21
+ ub = 2.069398670e-18 lub = -1.459027940e-24 wub = -2.553784995e-24 pub = 8.591000067e-30
+ uc = 1.754519487e-10 luc = -9.580631468e-16 wuc = -8.340638805e-16 puc = 6.314499858e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.662226723e+00 la0 = -3.288378617e-06 wa0 = -1.750769145e-06 pa0 = 1.661615534e-11
+ ags = 5.386641407e-01 lags = -8.129136481e-07 wags = -9.003366653e-07 pags = 6.831550788e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 1.461553941e-23 lb1 = -5.811337240e-29 wb1 = -7.243873489e-29 pb1 = 2.880262616e-34
+ keta = -2.849915097e-02 lketa = 1.056234113e-07 wketa = 8.996208595e-08 pketa = -3.590038095e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.019244331e+00 lpclm = 7.340044362e-06 wpclm = 3.396067243e-06 ppclm = -2.013478054e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 2.814622145e-03 lpdiblc2 = -3.119533207e-10 wpdiblc2 = 1.682108545e-09 ppdiblc2 = 3.114661224e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.004186824e+09 lpscbe1 = -8.013440292e+02 wpscbe1 = -2.049098704e+03 ppscbe1 = 8.074241626e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.596744755e-01 lkt1 = -2.008316174e-07 wkt1 = -3.565658870e-07 pkt1 = 1.280668045e-12
+ kt2 = -3.215028598e-02 lkt2 = -1.011128700e-07 wkt2 = -8.381152135e-08 pkt2 = 6.415196996e-13
+ at = 140000.0
+ ute = -1.119515970e+00 lute = -4.144964319e-06 wute = -4.551644711e-06 pute = 2.663844204e-11
+ ua1 = 1.919486860e-09 lua1 = -9.999862079e-15 wua1 = -9.374855506e-15 pua1 = 5.869887996e-20
+ ub1 = -2.193186578e-18 lub1 = 9.589233961e-24 wub1 = 9.024070989e-24 pub1 = -5.248415466e-29
+ uc1 = -2.774183419e-11 luc1 = 3.238684666e-16 wuc1 = 2.026400666e-16 puc1 = -1.451670441e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.080293429e-03 ltvoff = -5.288488554e-09 wtvoff = 1.824975995e-08 ptvoff = 5.356390680e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.12 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.423558564e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.201720421e-08 wvth0 = -3.553951225e-08 pvth0 = 1.497407486e-13
+ k1 = 5.755339035e-01 lk1 = -1.036218331e-07 wk1 = -1.766487394e-07 pk1 = 7.173232021e-13
+ k2 = -4.936388432e-02 lk2 = 4.110715310e-08 wk2 = 9.382282683e-08 pk2 = -3.374049164e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-8.431584123e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.558632845e-07 wvoff = -6.606846414e-07 pvoff = 1.290247154e-12
+ nfactor = 1.733761620e+00 lnfactor = 1.136590261e-06 wnfactor = 4.174084264e-06 pnfactor = -8.257074658e-12
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386683513e-01 letab = 2.730347037e-07 wetab = -1.176909134e-11 petab = 4.679550776e-17
+ u0 = 3.423494189e-02 lu0 = -7.424244779e-09 wu0 = -2.614048246e-09 pu0 = 6.477252463e-15
+ ua = -4.089115672e-10 lua = -1.590447614e-15 wua = -1.212818208e-15 pua = 6.355166684e-21
+ ub = 1.219303835e-18 lub = 1.921064737e-24 wub = 2.118126316e-24 pub = -9.985154686e-30
+ uc = -2.097160150e-10 luc = 5.734170597e-16 wuc = 1.541281884e-15 puc = -3.130197947e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 3.993356874e-01 la0 = 1.733047892e-06 wa0 = 5.675721869e-06 pa0 = -1.291258294e-11
+ ags = 2.441464682e-02 lags = 1.231812277e-06 wags = 1.668682765e-06 pags = -3.383219854e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.528191736e-05 lketa = -7.632325869e-09 wketa = -2.642739693e-08 pketa = 1.037766034e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.347779938e-01 lpclm = -3.180054735e-08 wpclm = -1.531916169e-06 ppclm = -5.404482921e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 1.329904060e-03 lpdiblc2 = 5.591487706e-09 wpdiblc2 = 4.126490088e-10 ppdiblc2 = 8.162204988e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.052652765e+08 lpscbe1 = -1.040490249e+01 wpscbe1 = -3.662674833e+01 ppscbe1 = 7.237943593e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.046813117e-01 lkt1 = -2.187831584e-08 wkt1 = -1.199379323e-08 pkt1 = -8.939746185e-14
+ kt2 = -5.814765051e-02 lkt2 = 2.256187043e-09 wkt2 = 8.157323401e-08 pkt2 = -1.607258004e-14
+ at = 1.677727274e+05 lat = -1.104281413e-01 wat = -2.095053599e-02 pat = 8.330218036e-8
+ ute = -2.533689068e+00 lute = 1.477980245e-06 wute = 3.783099279e-06 pute = -6.501633589e-12
+ ua1 = -1.721514169e-09 lua1 = 4.477253188e-15 wua1 = 1.111578179e-14 pua1 = -2.277468066e-20
+ ub1 = 1.239867144e-18 lub1 = -4.061054535e-24 wub1 = -1.001904353e-23 pub1 = 2.323385853e-29
+ uc1 = 6.727091944e-11 luc1 = -5.391516357e-17 wuc1 = -2.985607600e-16 puc1 = 5.411722084e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -7.829256732e-03 ltvoff = 9.617899398e-09 wtvoff = 4.066155142e-08 ptvoff = -8.375594021e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.13 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.276929598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.099308193e-08 wvth0 = 7.816108328e-08 pvth0 = -7.494709146e-14
+ k1 = 4.340894578e-01 lk1 = 1.758916280e-07 wk1 = 5.763314291e-07 pk1 = -7.706680160e-13
+ k2 = 7.716832658e-03 lk2 = -7.169210662e-08 wk2 = -2.556981581e-07 pk2 = 3.532960848e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.133108041e+00 ldsub = -1.725380231e-06 wdsub = -6.073585748e-06 pdsub = 1.200223145e-11
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.825196526e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.820080249e-08 wvoff = 1.965840146e-07 pvoff = -4.038322989e-13
+ nfactor = 2.768652783e+00 lnfactor = -9.084954210e-07 wnfactor = -1.727731173e-06 pnfactor = 3.405715291e-12
+ eta0 = -6.411041806e-03 leta0 = 1.365715851e-08 weta0 = 3.428240498e-08 peta0 = -6.774669465e-14
+ etab = -9.632053257e-04 letab = 9.106073408e-10 wetab = 1.939510043e-09 petab = -3.809197436e-15
+ u0 = 3.437662893e-02 lu0 = -7.704237635e-09 wu0 = 2.500804540e-09 pu0 = -3.630392263e-15
+ ua = -9.299748179e-10 lua = -5.607557664e-16 wua = 3.545575809e-15 pua = -3.048067035e-21
+ ub = 2.074615850e-18 lub = 2.308518719e-25 wub = -5.362545924e-24 pub = 4.797671032e-30
+ uc = 7.461009665e-11 luc = 1.154999470e-17 wuc = 8.920838520e-17 puc = -2.607032319e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.043538777e+04 lvsat = 1.177077746e-01 wvsat = 2.765056110e-01 pvsat = -5.464126921e-7
+ a0 = 2.487155610e+00 la0 = -2.392768220e-06 wa0 = -8.313672507e-06 pa0 = 1.473236291e-11
+ ags = 1.216823438e+00 lags = -1.124549661e-06 wags = -6.166359258e-06 pags = 1.209988875e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.144506780e-02 lketa = -1.093249755e-07 wketa = 8.223904274e-08 pketa = -1.109630600e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.096795738e+00 lpclm = -5.495832446e-07 wpclm = -2.602847633e-06 ppclm = 1.575857928e-12
+ pdiblc1 = -1.884416637e-01 lpdiblc1 = 1.143079395e-06 wpdiblc1 = 1.870182013e-06 ppdiblc1 = -3.695734003e-12
+ pdiblc2 = 6.815002987e-03 lpdiblc2 = -5.247813747e-09 wpdiblc2 = -8.490490509e-09 ppdiblc2 = 2.575601950e-14
+ pdiblcb = -4.898724213e-02 lpdiblcb = 4.740205271e-08 wpdiblcb = -1.593947540e-09 ppdiblcb = 3.149857116e-15
+ drout = 8.528408000e-01 ldrout = -5.786932471e-7
+ pscbe1 = 2.326916344e+09 lpscbe1 = -3.017394357e+03 wpscbe1 = -6.962207507e+03 ppscbe1 = 1.375826889e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.850882118e-07 lalpha0 = -7.017025985e-13 walpha0 = -2.019271745e-11 palpha0 = 3.990355590e-17
+ alpha1 = 8.168113760e-01 lalpha1 = 6.558523468e-8
+ beta0 = 1.182421474e+01 lbeta0 = 4.022988540e-06 wbeta0 = -4.661152279e-06 pbeta0 = 9.211070820e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.599484662e-01 lkt1 = 8.733709777e-08 wkt1 = -9.806652819e-08 pkt1 = 8.069396833e-14
+ kt2 = -8.698809060e-02 lkt2 = 5.924881895e-08 wkt2 = 1.457790957e-07 pkt2 = -1.429520948e-13
+ at = 1.562147447e+05 lat = -8.758799562e-02 wat = 6.308299700e-02 pat = -8.275950939e-8
+ ute = -2.561971268e+00 lute = 1.533869719e-06 wute = 2.695685041e-07 pute = 4.415810628e-13
+ ua1 = -8.561527015e-10 lua1 = 2.767181240e-15 wua1 = -2.339774547e-15 pua1 = 3.815328618e-21
+ ub1 = -3.464362798e-19 lub1 = -9.263032314e-25 wub1 = 4.605306503e-24 pub1 = -5.665846047e-30
+ uc1 = 1.177503932e-11 luc1 = 5.575224298e-17 wuc1 = 3.960554356e-17 puc1 = -1.270903981e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.504134558e-04 ltvoff = -4.766084838e-09 wtvoff = -1.936384505e-08 ptvoff = 3.486240667e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.14 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.616193217e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.876338769e-09 wvth0 = -6.290182826e-08 pvth0 = 6.274949477e-14
+ k1 = 7.174267341e-01 lk1 = -1.006840875e-07 wk1 = -2.822257427e-07 pk1 = 6.740054740e-14
+ k2 = -1.119025819e-01 lk2 = 4.507271025e-08 wk2 = 1.721231264e-07 pk2 = -6.431567268e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.707103633e+00 ldsub = 1.047052631e-06 wdsub = 1.278612866e-05 pdsub = -6.407414734e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.502744019e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 6.725052428e-09 wvoff = -3.651045665e-08 pvoff = -1.763003941e-13
+ nfactor = 1.471687587e+00 lnfactor = 3.575189979e-07 wnfactor = 3.607565500e-06 pnfactor = -1.802259862e-12
+ eta0 = -4.518150604e-01 leta0 = 4.484320556e-07 weta0 = -6.856480996e-08 peta0 = 3.264617435e-14
+ etab = 2.383608940e-04 letab = -2.622847026e-10 wetab = -3.831943721e-09 petab = 1.824526356e-15
+ u0 = 2.977408126e-02 lu0 = -3.211525165e-09 wu0 = -8.780563453e-09 pu0 = 7.381757165e-15
+ ua = -1.278540520e-09 lua = -2.205082364e-16 wua = -6.451937388e-17 pua = 4.758768363e-22
+ ub = 2.255126144e-18 lub = 5.464927589e-26 wub = -1.969794008e-25 pub = -2.446244123e-31
+ uc = 8.709476103e-11 luc = -6.367356515e-19 wuc = -3.273185511e-16 puc = 1.458837056e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.818354983e+05 lvsat = -3.984068376e-02 wvsat = -6.775515871e-01 pvsat = 3.848768850e-7
+ a0 = -1.358340181e+00 la0 = 1.360958660e-06 wa0 = 1.323417577e-05 pa0 = -6.301267513e-12
+ ags = -1.063868996e+00 lags = 1.101716328e-06 wags = 1.216136698e-05 pags = -5.790464627e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.110229117e-02 lketa = 2.005927328e-08 wketa = -1.416725565e-07 pketa = 1.076051128e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.650604639e-01 lpclm = 2.623034991e-07 wpclm = -7.918838127e-08 ppclm = -8.875767193e-13
+ pdiblc1 = 6.792427227e-01 lpdiblc1 = 2.961014293e-07 wpdiblc1 = -1.745617576e-06 ppdiblc1 = -1.662218555e-13
+ pdiblc2 = -1.452074582e-03 lpdiblc2 = 2.821978283e-09 wpdiblc2 = 4.188817168e-08 ppdiblc2 = -2.342040629e-14
+ pdiblcb = 2.297448426e-02 lpdiblcb = -2.284237904e-08 wpdiblcb = 3.187895080e-09 ppdiblcb = -1.517871612e-15
+ drout = 1.020293091e+00 ldrout = -7.421494565e-07 wdrout = -6.870374051e-06 pdrout = 6.706419445e-12
+ pscbe1 = -1.461636461e+09 lpscbe1 = 6.807484247e+02 wpscbe1 = 9.998067113e+03 ppscbe1 = -2.797265733e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.045363005e-05 lalpha0 = 1.963972049e-11 walpha0 = 1.383882472e-10 palpha0 = -1.148930326e-16
+ alpha1 = 9.163772480e-01 lalpha1 = -3.160459735e-8
+ beta0 = 1.569617265e+00 lbeta0 = 1.403287030e-05 wbeta0 = 9.041675896e-05 pbeta0 = -8.359790114e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.686553668e-01 lkt1 = -1.777383129e-09 wkt1 = -1.171499994e-09 pkt1 = -1.388875692e-14
+ kt2 = -1.757666685e-02 lkt2 = -8.506170576e-09 wkt2 = 2.911051178e-09 pkt2 = -3.493453254e-15
+ at = 7.989657716e+04 lat = -1.309108480e-02 wat = -4.915933551e-02 pat = 2.680427210e-8
+ ute = -6.803264328e-01 lute = -3.028715436e-07 wute = 2.142545094e-06 pute = -1.386698813e-12
+ ua1 = 2.582253735e-09 lua1 = -5.891710656e-16 wua1 = 4.534728970e-15 pua1 = -2.895121747e-21
+ ub1 = -1.239485765e-18 lub1 = -5.456547926e-26 wub1 = -3.366333665e-24 pub1 = 2.115558900e-30
+ uc1 = 1.498316505e-10 luc1 = -7.900978524e-17 wuc1 = -1.926657220e-16 puc1 = 9.963794597e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.441073950e-03 ltvoff = 9.840009341e-10 wtvoff = 2.011994366e-08 ptvoff = -3.679140905e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.15 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.190770893e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.948137287e-08 wvth0 = 5.867510028e-08 pvth0 = 4.862342318e-15
+ k1 = 2.822878334e-01 lk1 = 1.065012081e-07 wk1 = -3.214225439e-07 pk1 = 8.606355554e-14
+ k2 = 4.626208449e-02 lk2 = -3.023518136e-08 wk2 = 9.109183317e-08 pk2 = -2.573375684e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.873282620e-01 ldsub = 4.981820621e-08 wdsub = -9.651936128e-07 pdsub = 1.400848462e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.158305598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.674900752e-09 wvoff = -4.237090346e-07 pvoff = 8.058787995e-15
+ nfactor = 2.212878512e+00 lnfactor = 4.611315425e-09 wnfactor = -1.472278410e-06 pnfactor = 6.164366981e-13
+ eta0 = 0.49
+ etab = -2.569930338e-04 letab = -2.642886484e-11 wetab = 3.246611503e-09 petab = -1.545828615e-15
+ u0 = 2.669426170e-02 lu0 = -1.745112198e-09 wu0 = 1.892265732e-08 pu0 = -5.808743560e-15
+ ua = -1.349419498e-09 lua = -1.867602034e-16 wua = 1.518287228e-15 pua = -2.777543679e-22
+ ub = 1.999102462e-18 lub = 1.765513675e-25 wub = -2.100701032e-25 pub = -2.383914576e-31
+ uc = 4.031218941e-12 luc = 3.891280702e-17 wuc = 5.360116115e-16 puc = -2.651788647e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.247011095e+04 lvsat = 2.175483432e-02 wvsat = 2.935587506e-01 pvsat = -7.750370670e-8
+ a0 = 1.5
+ ags = 2.363013912e+00 lags = -5.299459918e-07 wags = -3.898278820e-12 pags = 1.856110885e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.540973132e-02 lketa = -6.457959399e-09 wketa = 6.363471476e-08 pketa = 9.850929874e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.211362672e+00 lpclm = -1.882650489e-07 wpclm = -3.909760516e-06 ppclm = 9.362965747e-13
+ pdiblc1 = 3.226103049e+00 lpdiblc1 = -9.165504588e-07 wpdiblc1 = -9.936612421e-06 ppdiblc1 = 3.733805666e-12
+ pdiblc2 = 6.207590322e-03 lpdiblc2 = -8.250639262e-10 wpdiblc2 = -1.378271132e-08 ppdiblc2 = 3.086505259e-15
+ pdiblcb = 6.042263145e-01 lpdiblcb = -2.995973005e-07 wpdiblcb = -3.118623057e-06 ppdiblcb = 1.484888708e-12
+ drout = -1.929948742e+00 ldrout = 6.625668886e-07 wdrout = 1.374074810e-05 pdrout = -3.107277813e-12
+ pscbe1 = -7.843924541e+08 lpscbe1 = 3.582881720e+02 wpscbe1 = 7.852695801e+03 ppscbe1 = -1.775777218e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.138540030e-05 lalpha0 = -9.804068065e-12 walpha0 = -2.250088190e-10 palpha0 = 5.813339291e-17
+ alpha1 = 0.85
+ beta0 = 4.244059302e+01 lbeta0 = -5.427272610e-06 wbeta0 = -1.665082017e-04 pbeta0 = 3.873332194e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.143827816e-01 lkt1 = -2.761851474e-08 wkt1 = -3.400134792e-07 pkt1 = 1.474461077e-13
+ kt2 = -1.068137071e-03 lkt2 = -1.636647591e-08 wkt2 = -2.191664868e-07 pkt2 = 1.022456574e-13
+ at = 7.917893229e+04 lat = -1.274938825e-02 wat = -6.070965093e-03 pat = 6.288347764e-9
+ ute = -1.212504931e+00 lute = -4.948220236e-08 wute = -5.005194258e-06 pute = 2.016597211e-12
+ ua1 = 1.746611269e-09 lua1 = -1.912916045e-16 wua1 = -6.466229626e-15 pua1 = 2.342830675e-21
+ ub1 = -2.103656553e-18 lub1 = 3.568973429e-25 wub1 = 3.572949936e-24 pub1 = -1.188483836e-30
+ uc1 = -1.358491248e-10 luc1 = 5.701311637e-17 wuc1 = 1.965021153e-16 puc1 = -8.565887140e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.585236814e-03 ltvoff = -3.757659364e-10 wtvoff = 7.279881281e-09 ptvoff = 2.434475036e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.16 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.109627752e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.764643433e-08 wvth0 = 2.989672687e-07 pvth0 = -4.947636747e-14
+ k1 = 4.580806325e-01 lk1 = 6.674812771e-08 wk1 = 1.733198696e-07 pk1 = -2.581551488e-14
+ k2 = 1.519391041e-02 lk2 = -2.320954874e-08 wk2 = -1.126201484e-07 pk2 = 2.033285583e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.052696561e+00 ldsub = -1.006455195e-07 wdsub = -9.748341775e-07 pdsub = 1.422649249e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {1.511242929e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -7.004300334e-08 wvoff = -1.961287216e-06 pvoff = 3.557605676e-13
+ nfactor = 1.634009772e+00 lnfactor = 1.355143767e-07 wnfactor = 4.252274630e-06 pnfactor = -6.780908282e-13
+ eta0 = 1.550355063e+00 leta0 = -2.397844526e-07 weta0 = -2.539778355e-07 peta0 = 5.743353180e-14
+ etab = 7.951944849e-02 letab = -1.806675425e-08 wetab = -1.331586887e-07 petab = 2.930032036e-14
+ u0 = -1.388581463e-02 lu0 = 7.431503943e-09 wu0 = 2.628088808e-08 pu0 = -7.472704432e-15
+ ua = -5.194822301e-09 lua = 6.828238050e-16 wua = 8.593040434e-17 pua = 4.615307479e-23
+ ub = 4.384694130e-18 lub = -3.629167898e-25 wub = 2.765827803e-24 pub = -9.113491065e-31
+ uc = 3.482642912e-10 luc = -3.893068301e-17 wuc = -1.862306271e-15 puc = 2.771671479e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.102388178e+04 lvsat = 1.755915880e-02 wvsat = 3.008783691e-01 pvsat = -7.915893596e-8
+ a0 = 1.5
+ ags = -2.725049684e+00 lags = 6.206483575e-07 wags = 1.392242436e-11 pags = -2.173791649e-18
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.132303484e-01 lketa = 1.340144366e-08 wketa = 5.300964428e-07 pketa = -9.563285946e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.175664524e+00 lpclm = -1.801924126e-07 wpclm = -3.364135541e-06 ppclm = 8.129111254e-13
+ pdiblc1 = -3.504829723e+00 lpdiblc1 = 6.055557544e-07 wpdiblc1 = 2.121927084e-05 ppdiblc1 = -3.311661150e-12
+ pdiblc2 = -8.867346784e-03 lpdiblc2 = 2.583922051e-09 wpdiblc2 = -1.823973298e-08 ppdiblc2 = 4.094398308e-15
+ pdiblcb = -2.245021456e+00 lpdiblcb = 3.447201932e-07 wpdiblcb = 1.190062844e-05 ppdiblcb = -1.911504749e-12
+ drout = 2.107148649e+00 ldrout = -2.503661669e-07 wdrout = -3.309056973e-06 pdrout = 7.482969076e-13
+ pscbe1 = 8.184696982e+08 lpscbe1 = -4.176663670e+00 wpscbe1 = -6.481001347e+01 ppscbe1 = 1.465587721e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.095849207e-06 lalpha0 = -1.145422138e-12 walpha0 = 3.763936372e-11 palpha0 = -1.260816547e-18
+ alpha1 = -2.783651019e+00 lalpha1 = 8.216993069e-07 walpha1 = 1.998416412e-05 palpha1 = -4.519138937e-12
+ beta0 = 4.486413993e+01 lbeta0 = -5.975323815e-06 wbeta0 = -1.149999148e-04 pbeta0 = 2.708544396e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.848447432e-01 lkt1 = 5.615627142e-08 wkt1 = 1.534668965e-06 pkt1 = -2.764870815e-13
+ kt2 = -1.553590431e-01 lkt2 = 1.852425241e-08 wkt2 = 7.440012128e-07 pkt2 = -1.155612335e-13
+ at = 3.846530241e+04 lat = -3.542570839e-03 wat = -2.430506920e-01 pat = 5.987799529e-8
+ ute = -6.059333123e-01 lute = -1.866498818e-07 wute = 1.299739770e-05 pute = -2.054436924e-12
+ ua1 = 4.223758656e-09 lua1 = -7.514638060e-16 wua1 = 1.204986547e-14 pua1 = -1.844325005e-21
+ ub1 = -4.489634735e-18 lub1 = 8.964529052e-25 wub1 = -2.407922044e-25 pub1 = -3.260594437e-31
+ uc1 = -9.851794355e-11 luc1 = 4.857119238e-17 wuc1 = 6.668615295e-16 puc1 = -1.920240679e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.831117902e-02 ltvoff = 2.954299729e-09 wtvoff = 8.315265643e-08 ptvoff = -1.472309084e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.17 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {7.253131642e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -3.550064667e-08 wvth0 = -6.814164349e-08 pvth0 = 7.842549637e-15
+ k1 = 8.024594106e-01 lk1 = 1.297820280e-08 wk1 = 1.181647507e-07 pk1 = -1.720381524e-14
+ k2 = -9.559405252e-02 lk2 = -5.911559364e-09 wk2 = -2.318175464e-07 pk2 = 3.894386077e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.439592925e+00 ldsub = -1.610539701e-07 wdsub = -5.121179048e-06 pdsub = 7.896586276e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 6.411402419e-02 lcdscd = -9.167371879e-09 wcdscd = -2.504924994e-07 pcdscd = 3.911089689e-14
+ cit = 0.0
+ voff = {3.133011516e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.133881960e-08 wvoff = -1.793968257e-06 pvoff = 3.296360546e-13
+ nfactor = 5.830433880e+00 lnfactor = -5.196984977e-07 wnfactor = -1.794551392e-05 pnfactor = 2.787783085e-12
+ eta0 = 7.206115648e-02 leta0 = -8.969555154e-09 weta0 = 5.975626641e-07 peta0 = -7.552259564e-14
+ etab = 3.506506218e-02 letab = -1.112582418e-08 wetab = -2.497332410e-08 petab = 1.240869027e-14
+ u0 = 7.460606954e-02 lu0 = -6.385264884e-09 wu0 = 8.413922277e-08 pu0 = -1.650647338e-14
+ ua = 6.033562110e-09 lua = -1.070331223e-15 wua = 4.584847861e-16 pua = -1.201607616e-23
+ ub = -5.149634739e-18 lub = 1.125735182e-24 wub = 6.867891660e-24 pub = -1.551828949e-30
+ uc = 1.721098632e-10 luc = -1.142663524e-17 wuc = 3.768785961e-16 puc = -7.245022046e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.843250382e+05 lvsat = -1.574483056e-02 wvsat = -1.257213226e+00 pvsat = 1.641152534e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.086656882e+00 lketa = 1.653883689e-07 wketa = 5.480040346e-06 pketa = -8.684973007e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -8.711599916e-01 lpclm = 1.393905800e-07 wpclm = 1.147277413e-05 ppclm = -1.503664604e-12
+ pdiblc1 = -1.280695971e-01 lpdiblc1 = 7.832193538e-08 wpdiblc1 = 3.152457680e-06 ppdiblc1 = -4.907812111e-13
+ pdiblc2 = -6.906294732e-03 lpdiblc2 = 2.277731228e-09 wpdiblc2 = 8.833404804e-08 ppdiblc2 = -1.254560557e-14
+ pdiblcb = -5.667230242e-01 lpdiblcb = 8.267738936e-08 wpdiblcb = 8.161113285e-07 ppdiblcb = -1.808125852e-13
+ drout = -2.487432580e-01 ldrout = 1.174733719e-07 wdrout = 1.199121755e-05 pdrout = -1.640626755e-12
+ pscbe1 = 8.143741681e+08 lpscbe1 = -3.537203979e+00 wpscbe1 = 2.825952501e+01 ppscbe1 = 1.243717468e-7
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.219442353e-05 lalpha0 = 2.803299886e-12 walpha0 = 1.538681049e-10 palpha0 = -1.940830728e-17
+ alpha1 = 9.328519045e+00 lalpha1 = -1.069446478e-06 walpha1 = -4.662971627e-05 palpha1 = 5.881685892e-12
+ beta0 = -2.395538075e+01 lbeta0 = 4.769880867e-06 wbeta0 = 3.043272422e-04 pbeta0 = -3.838662102e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.269357921e-01 lkt1 = 4.711459942e-08 wkt1 = 5.845589058e-07 pkt1 = -1.281406973e-13
+ kt2 = -6.472487730e-02 lkt2 = 4.372996302e-09 wkt2 = 1.930320397e-09 pkt2 = 3.027473130e-16
+ at = 2.162270652e+05 lat = -3.129758143e-02 wat = -1.159255683e+00 pat = 2.029305778e-7
+ ute = -9.375262849e+00 lute = 1.182558155e-06 wute = -8.358412305e-07 pute = 1.054296695e-13
+ ua1 = -1.321109607e-08 lua1 = 1.970744671e-15 wua1 = 1.372150595e-14 pua1 = -2.105328263e-21
+ ub1 = 8.031610843e-18 lub1 = -1.058564294e-24 wub1 = -6.900660490e-24 pub1 = 7.137857510e-31
+ uc1 = 2.439604408e-10 luc1 = -4.902012639e-18 wuc1 = -1.576303213e-15 puc1 = 1.582147024e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.687398671e-03 ltvoff = -9.488781963e-10 wtvoff = -3.690710632e-08 ptvoff = 4.022560272e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.18 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.363541752e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.771090359e-08 wvth0 = -3.596473666e-09 pvth0 = 3.595615404e-13
+ k1 = 5.438271891e-01 lk1 = -2.960832397e-07 wk1 = -1.658124366e-08 pk1 = 1.657728671e-12
+ k2 = -3.184284608e-02 lk2 = 9.431899429e-08 wk2 = 5.460897688e-09 pk2 = -5.459594500e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.797876101e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.658593950e-07 wvoff = 2.020996851e-08 pvoff = -2.020514560e-12
+ nfactor = 2.297782889e+00 lnfactor = 6.955451030e-07 wnfactor = -1.319499723e-07 pnfactor = 1.319184838e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.233087997e-02 lu0 = 1.021856337e-08 wu0 = 1.044550592e-09 pu0 = -1.044301320e-13
+ ua = -7.611659229e-10 lua = 2.501755769e-16 wua = -3.238132445e-17 pua = 3.237359697e-21
+ ub = 1.678526098e-18 lub = -4.333064184e-25 wub = 8.453359517e-26 pub = -8.451342208e-30
+ uc = 5.878403900e-11 luc = -9.539761888e-16 wuc = -4.424979731e-17 puc = 4.423923754e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.316726418e+00 la0 = -1.897888769e-06 wa0 = -1.179553725e-07 pa0 = 1.179272236e-11
+ ags = 4.357006798e-01 lags = -5.255425323e-07 wags = -2.290639080e-08 pags = 2.290092441e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.777924617e-25 lb0 = -7.776068493e-29 wb0 = -3.854958778e-30 pb0 = 3.854038830e-34
+ b1 = 2.633549380e-24 lb1 = -5.260814057e-29
+ keta = -9.250464793e-03 lketa = 4.557560051e-08 wketa = -9.678114294e-10 pketa = 9.675804709e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.614369198e-02 lpclm = 1.016988051e-06 wpclm = -1.216325199e-08 ppclm = 1.216034935e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.773573112e-03 lpdiblc2 = 2.998140236e-08 wpdiblc2 = 1.337521605e-09 ppdiblc2 = -1.337202419e-13
+ pdiblcb = -9.427960644e-01 lpdiblcb = 9.175770416e-05 wpdiblcb = 4.548856114e-06 ppdiblcb = -4.547770575e-10
+ drout = 0.56
+ pscbe1 = 8.062271626e+08 lpscbe1 = -5.154069996e+03 wpscbe1 = -1.810776562e+02 ppscbe1 = 1.810344439e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.072159914e-01 lkt1 = -5.812621098e-07 wkt1 = -1.474444443e-08 pkt1 = 1.474092582e-12
+ kt2 = -4.362268116e-02 lkt2 = -1.690252377e-07 wkt2 = -8.136593605e-09 pkt2 = 8.134651888e-13
+ at = 140000.0
+ ute = -1.761372561e+00 lute = -5.201502322e-06 wute = -1.708599392e-07 pute = 1.708191652e-11
+ ua1 = 4.317087131e-10 lua1 = -5.567542354e-15 wua1 = -1.313097049e-16 pua1 = 1.312783691e-20
+ ub1 = -6.481907438e-19 lub1 = 8.568698527e-25 wub1 = -1.329744002e-25 pub1 = 1.329426672e-29
+ uc1 = 1.484440068e-11 luc1 = 9.850771891e-17 wuc1 = 3.401823218e-18 puc1 = -3.401011407e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.150962748e-03 ltvoff = 1.276322824e-08 wtvoff = -7.256608209e-10 ptvoff = 7.254876492e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.19 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.349669748e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} wvth0 = 1.440308042e-8
+ k1 = 5.290053417e-01 wk1 = 6.640420812e-8
+ k2 = -2.712126257e-02 wk2 = -2.186968566e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.880904869e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} wvoff = -8.093644740e-8
+ nfactor = 2.332601690e+00 wnfactor = 5.284304124e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.284241851e-02 wu0 = -4.183193754e-9
+ ua = -7.486422008e-10 wua = 1.296800320e-16
+ ub = 1.656834896e-18 wub = -3.385383246e-25
+ uc = 1.102824735e-11 wuc = 1.772106370e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.221718616e+00 wa0 = 4.723851400e-7
+ ags = 4.093921618e-01 wags = 9.173502141e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.114886529e-24 wb0 = 1.543825604e-29
+ b1 = 0.0
+ keta = -6.968962479e-03 wketa = 3.875870406e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.705384049e-02 wpclm = 4.871113007e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 4.274434057e-03 wpdiblc2 = -5.356477769e-9
+ pdiblcb = 3.650569948e+00 wpdiblcb = -1.821716117e-5
+ drout = 0.56
+ pscbe1 = 5.482158036e+08 wpscbe1 = 7.251759048e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.363138165e-01 wkt1 = 5.904823407e-8
+ kt2 = -5.208403914e-02 wkt2 = 3.258525515e-8
+ at = 140000.0
+ ute = -2.021758369e+00 wute = 6.842562112e-7
+ ua1 = 1.529990390e-10 wua1 = 5.258662831e-16
+ ub1 = -6.052960693e-19 wub1 = 5.325330192e-25
+ uc1 = 1.977567061e-11 wuc1 = -1.362354849e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.512038972e-03 wtvoff = 2.906110855e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.20 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.317640336e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.554709460e-08 wvth0 = -8.805852583e-09 pvth0 = 1.851176060e-13
+ k1 = 5.143584298e-01 lk1 = 1.168257617e-07 wk1 = 1.004324218e-07 pk1 = -2.714136603e-13
+ k2 = -2.034204504e-02 lk2 = -5.407196102e-08 wk2 = -2.747211236e-08 pk2 = 4.468571725e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.005353381e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 9.926182602e-08 wvoff = -8.367090685e-08 pvoff = 2.181042043e-14
+ nfactor = 2.254092912e+00 lnfactor = 6.261966897e-07 wnfactor = 8.999044232e-07 pnfactor = -2.962927231e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.235149550e-02 lu0 = 3.915668706e-09 wu0 = -2.590538075e-09 pu0 = -1.270323829e-14
+ ua = -6.610039312e-10 lua = -6.990147567e-16 wua = -2.620612688e-16 pua = 3.124581892e-21
+ ub = 1.468911821e-18 lub = 1.498900005e-24 wub = 4.223971663e-25 pub = -6.069324963e-30
+ uc = -1.023161189e-10 luc = 9.040500801e-16 wuc = 5.426329932e-16 puc = -2.914658410e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.642080790e-01 la0 = 2.053939065e-06 wa0 = 1.708808093e-06 pa0 = -9.861877627e-12
+ ags = 2.535761891e-01 lags = 1.242809389e-06 wags = 5.126396173e-07 pags = -3.357192300e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.211189646e-24 lb0 = 2.469653475e-29 wb0 = 3.078440744e-29 pb0 = -1.224029907e-34
+ b1 = 0.0
+ keta = -9.975873028e-03 lketa = 2.398352748e-08 wketa = -1.844503110e-09 pketa = 4.562647714e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.557238492e-01 lpclm = 3.372132351e-06 wpclm = 1.074726238e-07 ppclm = -4.686896653e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 5.687552554e-03 lpdiblc2 = -1.127122532e-08 wpdiblc2 = -1.255694473e-08 ppdiblc2 = 5.743190375e-14
+ pdiblcb = 7.304211445e+00 lpdiblcb = -2.914194148e-05 wpdiblcb = -3.632563876e-05 ppdiblcb = 1.444356800e-10
+ drout = 0.56
+ pscbe1 = 3.005663900e+08 lpscbe1 = 1.975285403e+03 wpscbe1 = 1.438242589e+03 ppscbe1 = -5.687516851e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.574596798e-01 lkt1 = 1.686622815e-07 wkt1 = 1.280851606e-07 pkt1 = -5.506479151e-13
+ kt2 = -6.250017945e-02 lkt2 = 8.308055170e-08 wkt2 = 6.661110936e-08 pkt2 = -2.713948407e-13
+ at = 140000.0
+ ute = -2.363712447e+00 lute = 2.727472228e-06 wute = 1.614943892e-06 pute = -7.423291513e-12
+ ua1 = -4.847675260e-10 lua1 = 5.086912859e-15 wua1 = 2.541307231e-15 pua1 = -1.607543110e-20
+ ub1 = -1.851937603e-19 lub1 = -3.350793150e-24 wub1 = -9.281076705e-25 pub1 = 1.165026879e-29
+ uc1 = 2.776052890e-11 luc1 = -6.368831567e-17 wuc1 = -7.244529657e-17 puc1 = 4.691702624e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.258641363e-03 ltvoff = -2.021133789e-09 wtvoff = 4.264856610e-09 ptvoff = -1.083754093e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.21 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.210822990e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.801912398e-08 wvth0 = 6.989823710e-08 pvth0 = -1.278205583e-13
+ k1 = 5.393348269e-01 lk1 = 1.751620993e-08 wk1 = 2.764092559e-09 pk1 = 1.169288997e-13
+ k2 = -2.707715366e-02 lk2 = -2.729225315e-08 wk2 = -1.663649516e-08 pk2 = 1.601829622e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.294571546e+00 ldsub = -2.920756371e-06 wdsub = -2.171600641e-06 pdsub = 8.634579485e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.234135064e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.902285346e-07 wvoff = 2.872261282e-08 pvoff = -4.250814993e-13
+ nfactor = 2.704196237e+00 lnfactor = -1.163475347e-06 wnfactor = -6.356633602e-07 pnfactor = 3.142699113e-12
+ eta0 = 2.746614598e-01 leta0 = -7.740004382e-07 weta0 = -5.754741697e-07 peta0 = 2.288163563e-12
+ etab = -2.401757413e-01 letab = 6.766418914e-07 wetab = 5.030874809e-07 petab = -2.000344244e-12
+ u0 = 3.538043505e-02 lu0 = -8.127806897e-09 wu0 = -8.291435383e-09 pu0 = 9.964304725e-15
+ ua = -8.425297392e-10 lua = 2.275654349e-17 wua = 9.363157329e-16 pua = -1.640328046e-21
+ ub = 2.041556609e-18 lub = -7.780135537e-25 wub = -1.957190308e-24 pub = 3.392238460e-30
+ uc = 1.663509328e-10 luc = -1.642066562e-16 wuc = -3.226119606e-16 puc = 5.256731990e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.397832596e+00 la0 = -3.646346988e-06 wa0 = -4.229392387e-06 pa0 = 1.374921508e-11
+ ags = 6.049505850e-01 lags = -1.543029957e-07 wags = -1.208617056e-06 pags = 3.486758324e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.077719703e-24 lb0 = -1.223743211e-29 wb0 = -1.525404677e-29 pb0 = 6.065216449e-35
+ b1 = 0.0
+ keta = -1.066629930e-02 lketa = 2.672875624e-08 wketa = 2.636204881e-08 pketa = -6.652660941e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.023645232e-01 lpclm = -4.373573176e-07 wpclm = -3.800094678e-07 ppclm = 1.469605428e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 3.244423889e-04 lpdiblc2 = 1.005323008e-08 wpdiblc2 = 5.396000590e-09 ppdiblc2 = -1.395144844e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 7.825561225e+08 lpscbe1 = 5.882867629e+01 wpscbe1 = 7.592622305e+01 ppscbe1 = -2.707617044e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.953629437e-01 lkt1 = -7.824278632e-08 wkt1 = -5.817825285e-08 pkt1 = 1.899607487e-13
+ kt2 = -4.019094801e-02 lkt2 = -5.623986592e-09 wkt2 = -7.425247400e-09 pkt2 = 2.298378271e-14
+ at = 1.619829214e+05 lat = -8.740708497e-02 wat = 7.745375618e-03 pat = -3.079666683e-8
+ ute = -1.522233160e+00 lute = -6.183638592e-07 wute = -1.229961432e-06 pute = 3.888438961e-12
+ ua1 = 1.248403606e-09 lua1 = -1.804411272e-15 wua1 = -3.603968216e-15 pua1 = 8.359019832e-21
+ ub1 = -1.501811367e-18 lub1 = 1.884257516e-24 wub1 = 3.569488326e-24 pub1 = -6.232784567e-30
+ uc1 = 3.168071888e-12 luc1 = 3.409463800e-17 wuc1 = 1.915102945e-17 puc1 = 1.049708130e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.953098593e-03 ltvoff = -1.479144865e-08 wtvoff = -7.822560190e-09 ptvoff = 3.722367216e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.22 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.570975671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -3.151943894e-09 wvth0 = -6.757644263e-08 pvth0 = 1.438481054e-13
+ k1 = 4.322980265e-01 lk1 = 2.290354845e-07 wk1 = 5.852102679e-07 pk1 = -1.034063955e-12
+ k2 = -5.211285152e-03 lk2 = -7.050218309e-08 wk2 = -1.916227605e-07 pk2 = 3.473984882e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.489410334e+00 ldsub = 2.580770446e-06 wdsub = 6.924354866e-06 pdsub = -9.340265647e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.034098289e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.691505265e-08 wvoff = -1.955065805e-07 pvoff = 1.802588180e-14
+ nfactor = 1.670124830e+00 lnfactor = 8.799903886e-07 wnfactor = 3.716883148e-06 pnfactor = -5.458524734e-12
+ eta0 = -2.287746183e-01 leta0 = 2.208577195e-07 weta0 = 1.136378997e-06 peta0 = -1.094691106e-12
+ etab = 8.131145842e-02 letab = 4.133946247e-08 wetab = -4.058369249e-07 petab = -2.041860044e-13
+ u0 = 3.495217252e-02 lu0 = -7.281501884e-09 wu0 = -3.517517877e-10 pu0 = -5.725589857e-15
+ ua = -3.458116995e-10 lua = -9.588258568e-16 wua = 6.502986599e-16 pua = -1.075119411e-21
+ ub = 1.130976655e-18 lub = 1.021416273e-24 wub = -6.856039699e-25 pub = 8.794109197e-31
+ uc = 1.502659292e-10 luc = -1.324205014e-16 wuc = -2.857632557e-16 puc = 4.528551467e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.427304155e+04 lvsat = 3.107860877e-02 wvsat = 5.923383665e-02 pvsat = -1.170541170e-7
+ a0 = -9.487937003e-01 la0 = 2.967041715e-06 wa0 = 8.715861215e-06 pa0 = -1.183236659e-11
+ ags = -3.775707774e-01 lags = 1.787292839e-06 wags = 1.735908092e-06 pags = -2.332023824e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -6.155439406e-24 lb0 = 6.008546000e-30 wb0 = 3.050809353e-29 pb0 = -2.978004839e-35
+ b1 = 0.0
+ keta = 9.343023049e-02 lketa = -1.789801438e-07 wketa = -1.258512634e-07 pketa = 2.342675965e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.227253434e+00 lpclm = -1.672222791e-06 wpclm = -3.249432765e-06 ppclm = 7.139976106e-12
+ pdiblc1 = 2.243127512e-01 lpdiblc1 = 3.274205370e-07 wpdiblc1 = -1.755452639e-07 ppdiblc1 = 3.469013155e-13
+ pdiblc2 = 3.212200966e-03 lpdiblc2 = 4.346626400e-09 wpdiblc2 = 9.366012297e-09 ppdiblc2 = -2.179673150e-14
+ pdiblcb = -4.944563519e-02 lpdiblcb = 4.830789974e-08 wpdiblcb = 6.779777293e-10 ppdiblcb = -1.339776198e-15
+ drout = 8.528408000e-01 ldrout = -5.786932471e-7
+ pscbe1 = 5.784538022e+08 lpscbe1 = 4.621626191e+02 wpscbe1 = 1.703665918e+03 ppscbe1 = -3.487396714e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -9.144845511e-06 lalpha0 = 1.813074251e-11 walpha0 = 2.704032152e-11 palpha0 = -5.343535280e-17
+ alpha1 = 1.086627438e+00 lalpha1 = -4.676079994e-07 walpha1 = -1.337284493e-06 palpha1 = 2.642656028e-12
+ beta0 = 7.449738725e+00 lbeta0 = 1.266754807e-05 wbeta0 = 1.701998445e-05 pbeta0 = -3.363380400e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.679801847e-01 lkt1 = 6.525875782e-08 wkt1 = -5.825906639e-08 pkt1 = 1.901204472e-13
+ kt2 = -7.282323658e-02 lkt2 = 5.886185362e-08 wkt2 = 7.557408473e-08 pkt2 = -1.410341855e-13
+ at = 1.771510203e+05 lat = -1.173813113e-01 wat = -4.068308861e-02 pat = 6.490456476e-8
+ ute = -3.275796075e+00 lute = 2.846914947e-06 wute = 3.807485547e-06 pute = -6.066241361e-12
+ ua1 = -2.531529433e-09 lua1 = 5.665250484e-15 wua1 = 5.963864993e-15 pua1 = -1.054831981e-20
+ ub1 = 5.443922638e-19 lub1 = -2.159319143e-24 wub1 = 1.901090271e-25 pub1 = 4.453285231e-31
+ uc1 = -1.039974794e-10 luc1 = 2.458683418e-16 wuc1 = 6.134067940e-16 puc1 = -1.069359396e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -8.108883971e-03 ltvoff = 5.092397326e-09 wtvoff = 1.809806632e-08 ptvoff = -1.399901103e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.23 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.091172689e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.368335253e-08 wvth0 = 1.973131510e-07 pvth0 = -1.147201630e-13
+ k1 = 9.874452943e-01 lk1 = -3.128637488e-07 wk1 = -1.620513872e-06 pk1 = 1.119022784e-12
+ k2 = -1.898654730e-01 lk2 = 1.097454172e-07 wk2 = 5.585292002e-07 pk2 = -3.848518462e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.876654397e+00 ldsub = -7.049665158e-07 wdsub = -4.975986760e-06 pdsub = 2.276086227e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-9.239979068e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.766234735e-08 wvoff = -3.233533504e-07 pvoff = 1.428217164e-13
+ nfactor = 3.284871242e+00 lnfactor = -6.962217151e-07 wnfactor = -5.379084013e-06 pnfactor = 3.420376267e-12
+ eta0 = -4.715281226e-01 leta0 = 4.578181542e-07 weta0 = 2.913868551e-08 peta0 = -1.387397716e-14
+ etab = 2.412787209e-01 letab = -1.148103413e-07 wetab = -1.198495941e-06 petab = 5.695569972e-13
+ u0 = 2.838838065e-02 lu0 = -8.743483456e-10 wu0 = -1.912640458e-09 pu0 = -4.201950233e-15
+ ua = -1.172891700e-09 lua = -1.514832936e-16 wua = -5.881447193e-16 pua = 1.337697550e-22
+ ub = 2.093119325e-18 lub = 8.223417673e-26 wub = 6.059720805e-25 pub = -3.813429598e-31
+ uc = -5.719003815e-11 luc = 7.008473667e-17 wuc = 3.877976020e-16 puc = -2.046318547e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.689074767e+04 lvsat = 1.876201159e-02 wvsat = -1.574158084e-01 pvsat = 9.442540093e-8
+ a0 = 2.653372056e+00 la0 = -5.491619571e-07 wa0 = -6.649001382e-06 pa0 = 3.165828922e-12
+ ags = 1.554786768e+00 lags = -9.895092559e-08 wags = -8.174294508e-07 pags = 1.603808716e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.738030033e-01 lketa = 8.187583615e-08 wketa = 3.177783144e-07 pketa = -1.987752051e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.385751826e+00 lpclm = 8.784257117e-07 wpclm = 8.102702856e-06 ppclm = -3.941252151e-12
+ pdiblc1 = -2.765528811e-01 lpdiblc1 = 8.163335119e-07 wpdiblc1 = 2.991574971e-06 ppdiblc1 = -2.744638762e-12
+ pdiblc2 = 9.419806541e-03 lpdiblc2 = -1.712840875e-09 wpdiblc2 = -1.199593703e-08 ppdiblc2 = -9.445637253e-16
+ pdiblcb = 2.389127038e-02 lpdiblcb = -2.327889391e-08 wpdiblcb = -1.355955459e-09 ppdiblcb = 6.456192082e-16
+ drout = -2.494552533e-01 ldrout = 4.972976131e-07 wdrout = -5.771431887e-07 pdrout = 5.633702437e-13
+ pscbe1 = 1.291806799e+09 lpscbe1 = -2.341669223e+02 wpscbe1 = -3.648774159e+03 ppscbe1 = 1.737312733e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.289806226e-05 lalpha0 = -1.314749331e-11 walpha0 = -7.647496508e-11 palpha0 = 4.760964499e-17
+ alpha1 = 3.767451235e-01 lalpha1 = 2.253336839e-07 walpha1 = 2.674568986e-06 palpha1 = -1.273458578e-12
+ beta0 = 3.253329128e+01 lbeta0 = -1.181741058e-05 wbeta0 = -6.304794120e-05 pbeta0 = 4.452338067e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.236107223e-01 lkt1 = 2.194812831e-08 wkt1 = 2.712027395e-07 pkt1 = -1.314790822e-13
+ kt2 = 9.325787446e-03 lkt2 = -2.132676610e-08 wkt2 = -1.304250988e-07 pkt2 = 6.004903355e-14
+ at = 4.960931399e+04 lat = 7.116739710e-03 wat = 1.009528817e-01 pat = -7.335140480e-8
+ ute = 1.007947713e+00 lute = -1.334601580e-06 wute = -6.225017667e-06 pute = 3.726846196e-12
+ ua1 = 5.416821995e-09 lua1 = -2.093421486e-15 wua1 = -9.514190675e-15 pua1 = 4.560367534e-21
+ ub1 = -1.388221491e-18 lub1 = -2.728252830e-25 wub1 = -2.629157462e-24 pub1 = 3.197316037e-30
+ uc1 = 3.920554572e-10 luc1 = -2.383467875e-16 wuc1 = -1.393195215e-15 puc1 = 8.893570623e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.577905663e-03 ltvoff = 6.695462834e-10 wtvoff = 5.929274217e-09 ptvoff = -2.120614980e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.24 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.476887610e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.229552344e-08 wvth0 = -8.313241307e-08 pvth0 = 1.881006612e-14
+ k1 = -4.462581406e-02 lk1 = 1.785424604e-07 wk1 = 1.298853683e-06 pk1 = -2.709932064e-13
+ k2 = 1.558766633e-01 lk2 = -5.487486060e-08 wk2 = -4.521889309e-07 pk2 = 9.638744188e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.153734590e-01 ldsub = 3.841554494e-08 wdsub = -6.085653180e-07 pdsub = 1.965996510e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.111653539e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.113787120e-09 wvoff = 4.879708947e-08 pvoff = -3.437250540e-14
+ nfactor = 1.287537738e+00 lnfactor = 2.547806702e-07 wnfactor = 3.113971414e-06 pnfactor = -6.234731718e-13
+ eta0 = 0.49
+ etab = 1.910278903e-03 letab = -8.384087608e-10 wetab = -7.494999385e-09 petab = 2.478572728e-15
+ u0 = 3.375043898e-02 lu0 = -3.427417349e-09 wu0 = -1.604974710e-08 pu0 = 2.529235177e-15
+ ua = -8.915624399e-10 lua = -2.854342821e-16 wua = -7.509814663e-16 pua = 2.113021923e-22
+ ub = 1.924065949e-18 lub = 1.627265745e-25 wub = 1.618320143e-25 pub = -1.698718852e-31
+ uc = 1.640827545e-10 luc = -3.527120574e-17 wuc = -2.572489332e-16 puc = 1.024980224e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.183893099e+05 lvsat = -9.969478556e-04 wvsat = -3.315538882e-02 pvsat = 3.526054178e-8
+ a0 = 1.5
+ ags = 2.547688899e+00 lags = -5.717073745e-07 wags = -9.153052131e-07 pags = 2.069830455e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.560495070e-02 lketa = -8.308109442e-09 wketa = -1.396456155e-07 pketa = 1.902079523e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.506056264e-01 lpclm = 5.168341970e-08 wpclm = 3.563941332e-07 ppclm = -2.529557012e-13
+ pdiblc1 = 1.826620147e+00 lpdiblc1 = -1.850628808e-07 wpdiblc1 = -3.000380505e-06 ppdiblc1 = 1.083469502e-13
+ pdiblc2 = 8.864730888e-03 lpdiblc2 = -1.448549374e-09 wpdiblc2 = -2.695224928e-08 ppdiblc2 = 6.176674961e-15
+ pdiblcb = -2.924087145e-01 lpdiblcb = 1.273229157e-07 wpdiblcb = 1.325352999e-06 ppdiblcb = -6.310482753e-13
+ drout = 6.095479465e-01 ldrout = 8.829526556e-08 wdrout = 1.154286377e-06 pdrout = -2.610257043e-13
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.465450645e-05 lalpha0 = 4.732636541e-12 walpha0 = 5.274076208e-11 palpha0 = -1.391461447e-17
+ alpha1 = 0.85
+ beta0 = -3.230690459e+00 lbeta0 = 5.211108629e-06 wbeta0 = 5.985155848e-05 pbeta0 = -1.399349550e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.446665968e-01 lkt1 = -1.564001184e-08 wkt1 = -1.899183510e-07 pkt1 = 8.807726938e-14
+ kt2 = -3.116452394e-02 lkt2 = -2.047871194e-09 wkt2 = -7.000030631e-08 pkt2 = 3.127861454e-14
+ at = 9.235246539e+04 lat = -1.323481343e-02 wat = -7.136271010e-02 pat = 8.694251837e-9
+ ute = -2.354879333e+00 lute = 2.665614384e-07 wute = 6.567354300e-07 pute = 4.501958030e-13
+ ua1 = 1.356030169e-09 lua1 = -1.599323086e-16 wua1 = -4.530399546e-15 pua1 = 2.187405161e-21
+ ub1 = -3.727401675e-18 lub1 = 8.409426132e-25 wub1 = 1.162068866e-23 pub1 = -3.587548696e-30
+ uc1 = -3.170077008e-10 luc1 = 9.926370828e-17 wuc1 = 1.094375105e-15 puc1 = -2.950647196e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.990807394e-03 ltvoff = -8.612833775e-11 wtvoff = -6.225605532e-10 ptvoff = 9.989494198e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.25 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.889840953e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -3.163388516e-08 wvth0 = -8.772839592e-08 pvth0 = 1.984938330e-14
+ k1 = 4.931050082e-01 lk1 = 5.694216317e-08 wk1 = -2.708135376e-10 pk1 = 2.278561067e-14
+ k2 = -1.765604210e-03 lk2 = -1.922626879e-08 wk2 = -2.856401140e-08 pk2 = 5.905970865e-16
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.949779736e-01 ldsub = -9.265390157e-08 wdsub = -1.931363806e-07 pdsub = 1.026562128e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -5.638404937e-03 lcdscd = 2.496180739e-09 wcdscd = 5.470944770e-08 pcdscd = -1.237177566e-14
+ cit = 0.0
+ voff = {-2.801629498e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.448905321e-08 wvoff = 1.762939818e-07 pvoff = -6.320414264e-14
+ nfactor = 2.273383696e+00 lnfactor = 3.184540849e-08 wnfactor = 1.083357161e-06 pnfactor = -1.642781871e-13
+ eta0 = 1.377471867e+00 leta0 = -2.006893380e-07 weta0 = 6.028800406e-07 peta0 = -1.363328809e-13
+ etab = -3.521303131e-02 letab = 7.556508117e-09 wetab = 4.354878357e-07 petab = -9.769579367e-14
+ u0 = -7.997993961e-03 lu0 = 6.013406282e-09 wu0 = -2.900811512e-09 pu0 = -4.442125222e-16
+ ua = -6.749666627e-09 lua = 1.039293966e-15 wua = 7.792177348e-15 pua = -1.720613569e-21
+ ub = 7.661363531e-18 lub = -1.134682951e-24 wub = -1.347426977e-23 pub = 2.913741628e-30
+ uc = -2.264736401e-10 luc = 5.304765511e-17 wuc = 9.862569928e-16 puc = -1.787034337e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.079762222e+04 lvsat = 5.242526038e-03 wvsat = 2.028741352e-01 pvsat = -1.811423068e-8
+ a0 = 1.5
+ ags = -2.725045681e+00 lags = 6.206477325e-07 wags = -5.916754457e-12 pags = 9.238183736e-19
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.781446191e-03 lketa = -6.538933426e-09 wketa = -6.967213643e-08 pketa = 3.197272573e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.388206768e-01 lpclm = 9.121221069e-09 wpclm = -2.077578437e-07 ppclm = -1.253806297e-13
+ pdiblc1 = 2.359042693e+00 lpdiblc1 = -3.054627857e-07 wpdiblc1 = -7.843734467e-06 ppdiblc1 = 1.203603642e-12
+ pdiblc2 = -1.570608770e-02 lpdiblc2 = 4.107797258e-09 wpdiblc2 = 1.565499552e-08 ppdiblc2 = -3.458356948e-15
+ pdiblcb = 1.120676856e+00 lpdiblcb = -1.922266030e-07 wpdiblcb = -4.780721519e-06 ppdiblcb = 7.497549918e-13
+ drout = 4.516027116e-01 ldrout = 1.240123692e-07 wdrout = 4.896295556e-06 pdrout = -1.107228692e-12
+ pscbe1 = 7.850767286e+08 lpscbe1 = 3.374688911e+00 wpscbe1 = 1.006949609e+02 ppscbe1 = -2.277075567e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.083252961e-05 lalpha0 = -1.030899845e-12 walpha0 = -7.058061165e-13 palpha0 = -1.828421326e-18
+ alpha1 = 1.837382488e+00 lalpha1 = -2.232827263e-07 walpha1 = -2.918981076e-06 palpha1 = 6.600867046e-13
+ beta0 = 9.327764020e+00 lbeta0 = 2.371189967e-06 wbeta0 = 6.112838551e-05 pbeta0 = -1.428223206e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.331906060e-01 lkt1 = 4.378453513e-09 wkt1 = 2.874000947e-07 pkt1 = -1.986161466e-14
+ kt2 = -2.650655854e-02 lkt2 = -3.101204857e-09 wkt2 = 1.053719629e-07 pkt2 = -8.379368922e-15
+ at = 1.150888746e+05 lat = -1.837633407e-02 wat = -6.228187239e-01 pat = 1.333983090e-7
+ ute = 1.987849026e+00 lute = -7.154857818e-07 wute = 1.418809837e-07 pute = 5.666229281e-13
+ ua1 = 5.008738400e-09 lua1 = -9.859411372e-16 wua1 = 8.159284493e-15 pua1 = -6.821892292e-22
+ ub1 = -2.016597456e-18 lub1 = 4.540681903e-25 wub1 = -1.249786236e-23 pub1 = 1.866523956e-30
+ uc1 = 3.321514218e-10 luc1 = -4.753453906e-17 wuc1 = -1.467657294e-15 puc1 = 2.843030389e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.570300860e-03 ltvoff = 2.710519966e-10 wtvoff = 1.009270736e-08 ptvoff = -1.424158405e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.26 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {7.573614292e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -4.231004857e-08 wvth0 = -2.269818826e-07 pvth0 = 4.159186570e-14
+ k1 = 7.069074261e-01 lk1 = 2.355990885e-08 wk1 = 5.917473316e-07 pk1 = -6.964973445e-14
+ k2 = -1.710019540e-01 lk2 = 7.197617925e-09 wk2 = 1.419252784e-07 pk2 = -2.602891866e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.289742177e-01 ldsub = -4.280339138e-09 wdsub = 3.833604585e-07 pdsub = 1.264430231e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 3.060418107e-02 lcdscd = -3.162591669e-09 wcdscd = -8.440829895e-08 pcdscd = 9.349512825e-15
+ cit = 0.0
+ voff = {-2.851824390e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.527277618e-08 wvoff = -2.252427817e-07 pvoff = -5.097985388e-16
+ nfactor = 3.347848293e+00 lnfactor = -1.359171958e-07 wnfactor = -5.641119659e-06 pnfactor = 8.856547257e-13
+ eta0 = 4.763329940e-01 leta0 = -5.998911901e-08 weta0 = -1.406122568e-06 peta0 = 1.773447504e-13
+ etab = 1.500326779e-01 letab = -2.136701594e-08 wetab = -5.947852485e-07 petab = 6.316692461e-14
+ u0 = 1.742846561e-01 lu0 = -2.244747756e-08 wu0 = -4.098959614e-07 pu0 = 6.310238219e-14
+ ua = 1.697280683e-08 lua = -2.664638150e-15 wua = -5.375949692e-14 pua = 7.889818645e-21
+ ub = -1.396242758e-17 lub = 2.241569298e-24 wub = 5.054657819e-23 pub = -7.082217490e-30
+ uc = 5.266491414e-10 luc = -6.454192351e-17 wuc = -1.380318047e-15 puc = 1.908041267e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -5.294991105e+04 lvsat = 2.768669089e-02 wvsat = 4.144165339e-01 pvsat = -5.114361464e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.519339594e-01 lketa = -9.150073022e-08 wketa = -2.641277947e-06 pketa = 4.047175174e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.605040018e+00 lpclm = -3.134900019e-07 wpclm = -5.756253401e-06 ppclm = 7.409392726e-13
+ pdiblc1 = 7.311991496e-01 lpdiblc1 = -5.129780627e-08 wpdiblc1 = -1.106320543e-06 ppdiblc1 = 1.516507813e-13
+ pdiblc2 = 1.462683294e-02 lpdiblc2 = -6.282636394e-10 wpdiblc2 = -1.839020505e-08 ppdiblc2 = 1.857324488e-15
+ pdiblcb = -8.436781848e-01 lpdiblcb = 1.144799357e-07 wpdiblcb = 2.188779206e-06 ppdiblcb = -3.384349734e-13
+ drout = 4.635200135e+00 ldrout = -5.291977980e-07 wdrout = -1.221498318e-05 pdrout = 1.564457925e-12
+ pscbe1 = 8.624336049e+08 lpscbe1 = -8.703504333e+00 wpscbe1 = -2.099365967e+02 ppscbe1 = 2.573001320e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.188879730e-05 lalpha0 = -2.757181256e-12 walpha0 = -6.462076899e-11 palpha0 = 8.151005317e-18
+ alpha1 = -1.453892472e+00 lalpha1 = 2.906037808e-07 walpha1 = 6.810955844e-06 palpha1 = -8.591067263e-13
+ beta0 = 6.931149233e+01 lbeta0 = -6.994429437e-06 wbeta0 = -1.579296821e-04 pbeta0 = 1.992061838e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.425863786e-01 lkt1 = 5.268627187e-08 wkt1 = 1.157755826e-06 pkt1 = -1.557554772e-13
+ kt2 = -1.167450682e-01 lkt2 = 1.098827508e-08 wkt2 = 2.597570561e-07 pkt2 = -3.248443984e-14
+ at = -2.489356391e+05 lat = 3.846099742e-02 wat = 1.146221855e+00 pat = -1.428126109e-7
+ ute = -2.170141203e+01 lute = 2.983260683e-06 wute = 6.025603010e-05 pute = -8.819359858e-12
+ ua1 = -2.584295612e-08 lua1 = 3.831119038e-15 wua1 = 7.632856654e-14 pua1 = -1.132586825e-20
+ ub1 = 1.540697490e-17 lub1 = -2.266378703e-24 wub1 = -4.345504462e-23 pub1 = 6.700054566e-30
+ uc1 = -4.011452666e-10 luc1 = 6.695947268e-17 wuc1 = 1.621022593e-15 puc1 = -1.979510838e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.125734085e-04 ltvoff = -2.219829368e-10 wtvoff = -1.717642506e-09 ptvoff = 4.198623815e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.27 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.307468172e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.816266804e-07 wvth0 = 1.298045784e-08 pvth0 = -2.592993912e-13
+ k1 = 5.344591002e-01 lk1 = 3.397603097e-07 wk1 = 1.111346905e-08 pk1 = -2.220041692e-13
+ k2 = -2.844478878e-02 lk2 = -1.213385104e-07 wk2 = -4.584717946e-09 pk2 = 9.158494921e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.167853073e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.971304284e-06 wvoff = -1.660426054e-07 pvoff = 3.316889666e-12
+ nfactor = 1.924376605e+00 lnfactor = 1.172546038e-05 wnfactor = 9.719443042e-07 pnfactor = -1.941569161e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.374692911e-02 lu0 = -4.633522903e-08 wu0 = -3.141689988e-09 pu0 = 6.275882647e-14
+ ua = -8.605860935e-10 lua = 3.112478025e-15 wua = 2.615327364e-16 pua = -5.224413510e-21
+ ub = 1.916544460e-18 lub = -7.475558700e-24 wub = -6.191158015e-25 pub = 1.236754145e-29
+ uc = 4.982766889e-11 luc = 4.223820340e-16 wuc = -1.777224155e-17 puc = 3.550207143e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.229676699e+00 la0 = 3.033020705e-06 wa0 = 1.393881458e-07 pa0 = -2.784436558e-12
+ ags = 4.341693491e-01 lags = 1.249177888e-07 wags = -1.837934537e-08 pags = 3.671483028e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.261963924e-25 lb0 = 5.260708209e-29
+ b1 = 7.785514628e-24 lb1 = -1.555244990e-28 wb1 = -1.523066213e-29 pb1 = 3.042497780e-34
+ keta = -1.595293910e-02 lketa = 2.056551011e-07 wketa = 1.884659271e-08 pketa = -3.764820991e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.115928690e-01 lpclm = 3.897820945e-06 wpclm = 3.654620441e-07 ppclm = -7.300519495e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.932071753e-03 lpdiblc2 = -9.379484098e-09 wpdiblc2 = 8.689549233e-10 ppdiblc2 = -1.735836173e-14
+ pdiblcb = 5.959123923e-01 lpdiblcb = -6.207642177e-05 wpdiblcb = -1.942890293e-22 ppdiblcb = 9.769962617e-27
+ drout = 0.56
+ pscbe1 = 8.920131824e+08 lpscbe1 = -1.967597506e+03 wpscbe1 = -4.346853224e+02 ppscbe1 = 8.683333118e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.844064645e-01 lkt1 = -6.379086479e-07 wkt1 = -8.217583833e-08 pkt1 = 1.641555722e-12
+ kt2 = -4.589540693e-02 lkt2 = 9.655954614e-08 wkt2 = -1.417775330e-09 pkt2 = 2.832167281e-14
+ at = 140000.0
+ ute = -1.647300853e+00 lute = -2.856570414e-06 wute = -5.080880770e-07 pute = 1.014963653e-11
+ ua1 = 6.731339193e-10 lua1 = -6.836910839e-15 wua1 = -8.450306964e-16 pua1 = 1.688044812e-20
+ ub1 = -1.039765919e-18 lub1 = 1.227745143e-23 wub1 = 1.024632243e-24 pub1 = -2.046819303e-29
+ uc1 = 1.306819906e-11 luc1 = 4.193256512e-17 wuc1 = 8.652776088e-18 puc1 = -1.728490319e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.079829591e-03 ltvoff = 9.090779106e-08 wtvoff = 7.932895507e-09 ptvoff = -1.584685995e-13
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.28 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.539839+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.55146741
+ k2 = -0.034518962
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.21546827+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.51135
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314274
+ ua = -7.0477628e-10
+ ub = 1.54232e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3815089
+ ags = 0.4404227
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -0.00052901
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.29 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.287853419e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 8.816548014e-8
+ k1 = 5.483309743e-01 lk1 = 2.501663785e-8
+ k2 = -2.963483658e-02 lk2 = -3.895644861e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.288380869e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.066394782e-7
+ nfactor = 2.558497033e+00 lnfactor = -3.760511442e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.147521304e-02 lu0 = -3.813632729e-10
+ ua = -7.496494897e-10 lua = 3.579148231e-16
+ ub = 1.611793036e-18 lub = -5.541263855e-25
+ uc = 8.123639508e-11 luc = -8.187021115e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.542234158e+00 la0 = -1.281966517e-6
+ ags = 4.269830621e-01 lags = 1.071963796e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.202027848e-24 lb0 = -1.670783420e-29
+ b1 = 0.0
+ keta = -1.059979967e-02 lketa = 3.941726389e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.193698668e-01 lpclm = 3.213592108e-06 wpclm = 1.110223025e-22 ppclm = -1.332267630e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.440006234e-03 lpdiblc2 = 8.155846848e-9
+ pdiblcb = -4.983398045e+00 lpdiblcb = 1.971526497e-5
+ drout = 0.56
+ pscbe1 = 7.870702449e+08 lpscbe1 = 5.141046490e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141332445e-01 lkt1 = -1.760138183e-8
+ kt2 = -3.996812420e-02 lkt2 = -8.722206193e-9
+ at = 140000.0
+ ute = -1.817437128e+00 lute = 2.164494252e-7
+ ua1 = 3.748619787e-10 lua1 = -3.508062434e-16
+ ub1 = -4.991379884e-19 lub1 = 5.900584965e-25
+ uc1 = 3.254985601e-12 luc1 = 9.501449495e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.840006479e-04 ltvoff = -5.687069897e-09 ptvoff = -3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.30 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.447262671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.478219384e-8
+ k1 = 5.402698164e-01 lk1 = 5.706889798e-8
+ k2 = -3.270465982e-02 lk2 = -2.675041390e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.136977172e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 4.643930903e-8
+ nfactor = 2.489175018e+00 lnfactor = -1.004173866e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.257575154e-02 lu0 = -4.757254045e-9
+ ua = -5.258090296e-10 lua = -5.321052884e-16
+ ub = 1.379512085e-18 lub = 3.694542658e-25
+ uc = 5.722333245e-11 luc = 1.360899167e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.671868096e-01 la0 = 1.004499947e-6
+ ags = 1.961204884e-01 lags = 1.025137370e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.082155696e-24 lb0 = 8.278934222e-30
+ b1 = 0.0
+ keta = -1.749000880e-03 lketa = 4.225284179e-09 pketa = -1.734723476e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.738214857e-01 lpclm = 5.975541666e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.149708243e-03 lpdiblc2 = 5.333975140e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.082391335e+08 lpscbe1 = -3.275991519e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.150424779e-01 lkt1 = -1.398614617e-8
+ kt2 = -4.270263241e-02 lkt2 = 2.150570337e-9
+ at = 1.646028932e+05 lat = -9.782444936e-2
+ ute = -1.938283263e+00 lute = 6.969500930e-7
+ ua1 = 2.931550244e-11 lua1 = 1.023133540e-15
+ ub1 = -2.943865257e-19 lub1 = -2.240611654e-25
+ uc1 = 9.646151264e-12 luc1 = 6.960235108e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.929819200e-04 ltvoff = -2.200067937e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.31 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.342389756e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.550650798e-8
+ k1 = 6.302528454e-01 lk1 = -1.207498050e-7
+ k2 = -7.003012197e-02 lk2 = 4.700977557e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.695424173e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.081756878e-8
+ nfactor = 2.927407845e+00 lnfactor = -9.664250529e-07 wnfactor = 3.552713679e-21
+ eta0 = 1.556200357e-01 leta0 = -1.494354750e-7
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 3.483318800e-02 lu0 = -9.218255501e-9
+ ua = -1.258399038e-10 lua = -1.322498677e-15
+ ub = 8.990623895e-19 lub = 1.318888206e-24
+ uc = 5.360287210e-11 luc = 2.076351371e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.430964044e+04 lvsat = -8.516435621e-3
+ a0 = 1.999457250e+00 la0 = -1.035406831e-6
+ ags = 2.096222212e-01 lags = 9.984561099e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.164311393e-24 lb0 = -4.064934266e-30
+ b1 = 0.0
+ keta = 5.085943942e-02 lketa = -9.973614859e-08 wketa = -1.994931997e-23 pketa = -4.423544864e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.280914582e-01 lpclm = 7.429649702e-7
+ pdiblc1 = 1.649323322e-01 lpdiblc1 = 4.447643207e-7
+ pdiblc2 = 6.380373791e-03 lpdiblc2 = -3.026395354e-9
+ pdiblcb = -4.921630060e-02 lpdiblcb = 4.785470340e-8
+ drout = 8.528408000e-01 ldrout = -5.786932471e-7
+ pscbe1 = 1.154740475e+09 lpscbe1 = -7.174936905e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.887283200e-09 lalpha0 = 5.555455173e-14
+ alpha1 = 6.342739440e-01 lalpha1 = 4.263040254e-7
+ beta0 = 1.320696502e+01 lbeta0 = 1.290485941e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.876870551e-01 lkt1 = 1.295694180e-7
+ kt2 = -4.725934087e-02 lkt2 = 1.115524596e-8
+ at = 1.633894479e+05 lat = -9.542651645e-2
+ ute = -1.987865646e+00 lute = 7.949316238e-7
+ ua1 = -5.141762198e-10 lua1 = 2.097147098e-15 pua1 = 8.271806126e-37
+ ub1 = 6.086990610e-19 lub1 = -2.008681104e-24 pub1 = -7.703719778e-46
+ uc1 = 1.034951732e-10 luc1 = -1.158560798e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.986982774e-03 ltvoff = 3.570537335e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.32 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.758609527e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.877797783e-9
+ k1 = 4.392858589e-01 lk1 = 6.565994532e-8
+ k2 = -9.358647387e-04 lk2 = -2.043561631e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.934635650e-01 ldsub = 6.494860950e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.017781756e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.351084606e-9
+ nfactor = 1.465327635e+00 lnfactor = 4.607640755e-7
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 1.977584763e-22 peta0 = -7.285838599e-29
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.774140568e-02 lu0 = -2.295711474e-9
+ ua = -1.371839134e-09 lua = -1.062339720e-16
+ ub = 2.298097091e-18 lub = -4.675993133e-26
+ uc = 7.398743477e-11 luc = 8.654082393e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.364284762e+04 lvsat = 5.070260485e-2
+ a0 = 4.042627414e-01 la0 = 5.217199554e-7
+ ags = 1.278280856e+00 lags = -4.470005522e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.631044528e-02 lketa = 1.463759397e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.355090508e+00 lpclm = -4.547529740e-7
+ pdiblc1 = 7.353854155e-01 lpdiblc1 = -1.120754702e-7
+ pdiblc2 = 5.362028211e-03 lpdiblc2 = -2.032351573e-9
+ pdiblcb = 2.343260119e-02 lpdiblcb = -2.306050500e-08 wpdiblcb = 3.903127821e-24 ppdiblcb = -2.385244779e-30
+ drout = -4.446812800e-01 ldrout = 6.878647659e-07 pdrout = 2.220446049e-28
+ pscbe1 = 5.756251585e+07 lpscbe1 = 3.535012140e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.970567686e-06 lalpha0 = 2.957074856e-12 walpha0 = -5.293955920e-28 palpha0 = -6.882142696e-34
+ alpha1 = 1.281452112e+00 lalpha1 = -2.054298828e-7
+ beta0 = 1.120652299e+01 lbeta0 = 3.243189417e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.318729451e-01 lkt1 = -2.252634408e-8
+ kt2 = -3.479216166e-02 lkt2 = -1.014416479e-9
+ at = 8.375791069e+04 lat = -1.769530623e-2
+ ute = -1.097743715e+00 lute = -7.394843689e-8
+ ua1 = 2.198525948e-09 lua1 = -5.508191447e-16
+ ub1 = -2.277567454e-18 lub1 = 8.087075466e-25
+ uc1 = -7.921055025e-11 luc1 = 6.248955431e-17 puc1 = -1.292469707e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.572253219e-03 ltvoff = -4.777871482e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.33 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.195681646e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.593277925e-8
+ k1 = 3.947279698e-01 lk1 = 8.687556041e-8
+ k2 = 2.918004145e-03 lk2 = -2.227058202e-08 pk2 = -1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.095184973e-01 ldsub = 1.049178783e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.946591176e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.274072440e-8
+ nfactor = 2.340878188e+00 lnfactor = 4.388293722e-8
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 2.832140781e-02 lu0 = -2.571871370e-9
+ ua = -1.145591476e-09 lua = -2.139586271e-16
+ ub = 1.978807687e-18 lub = 1.052652480e-25
+ uc = 7.706502979e-11 luc = -5.999455450e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.071740778e+05 lvsat = 1.093037903e-2
+ a0 = 1.5
+ ags = 2.238075265e+00 lags = -5.016927259e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.163195547e-02 lketa = -1.874083449e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.711604765e-01 lpclm = -3.388206463e-8
+ pdiblc1 = 8.117032664e-01 lpdiblc1 = -1.484131464e-7
+ pdiblc2 = -2.522103509e-04 lpdiblc2 = 6.407895190e-10
+ pdiblcb = 1.559088000e-01 lpdiblcb = -8.613719240e-08 ppdiblcb = 2.081668171e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.185727360e-06 lalpha0 = 2.584115772e-14
+ alpha1 = 0.85
+ beta0 = 1.701486070e+01 lbeta0 = 4.776307318e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.089088954e-01 lkt1 = 1.415324515e-8
+ kt2 = -5.484301818e-02 lkt2 = 8.532518139e-9
+ at = 6.821312074e+04 lat = -1.029387212e-2
+ ute = -2.132730218e+00 lute = 4.188458967e-7
+ ua1 = -1.764351194e-10 lua1 = 5.799853180e-16
+ ub1 = 2.034441167e-19 lub1 = -3.725913786e-25 pub1 = 1.925929944e-46
+ uc1 = 5.317860243e-11 luc1 = -5.456872969e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.201396422e-03 ltvoff = 2.517790134e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.34 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.221980462e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.086109844e-09 wvth0 = 4.053381990e-07 pvth0 = -9.166155898e-14
+ k1 = 4.930134021e-01 lk1 = 6.464968589e-8
+ k2 = -1.079110766e-02 lk2 = -1.917045832e-08 wk2 = -1.882078004e-09 pk2 = 4.256055914e-16
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.296255798e-01 ldsub = -5.792425694e-08 wdsub = 6.372491664e-11 pdsub = -1.441049775e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.286776183e-02 lcdscd = -1.688729789e-09 wcdscd = 1.387778781e-23
+ cit = 0.0
+ voff = {-2.123258593e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -8.745638097e-09 wvoff = -2.425158771e-08 pvoff = 5.484157039e-15
+ nfactor = 2.513344741e+00 lnfactor = 4.882040737e-09 wnfactor = 3.739646424e-07 pnfactor = -8.456686838e-14
+ eta0 = 1.581403705e+00 leta0 = -2.468056683e-07 weta0 = 1.573773112e-14 peta0 = -3.558867867e-21
+ etab = 1.433521275e-01 letab = -3.255841171e-08 wetab = -9.240112913e-08 petab = 2.089522174e-14
+ u0 = -8.777635972e-03 lu0 = 5.817557996e-09 wu0 = -5.959698682e-10 pu0 = 1.347702421e-16
+ ua = -4.117754007e-09 lua = 4.581543190e-16 wua = 1.150144447e-17 pua = -2.600890647e-24
+ ub = 2.543297387e-18 lub = -2.238619480e-26 wub = 1.656177044e-24 pub = -3.745212521e-31
+ uc = 2.061964889e-10 luc = -2.980121719e-17 wuc = -2.928379216e-16 puc = 6.622119624e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.362187155e+05 lvsat = -1.825125916e-02 wvsat = -2.270316253e-01 pvsat = 5.134002363e-8
+ a0 = 1.5
+ ags = -2.725047683e+00 lags = 6.206480450e-07 wags = -3.330669074e-22 pags = 4.163336342e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.859815628e-01 lketa = -7.369793403e-08 wketa = -8.921101337e-07 pketa = 2.017382172e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.289816123e-02 lpclm = 6.748618229e-08 wpclm = 1.317454603e-06 ppclm = -2.979239140e-13
+ pdiblc1 = -2.942002886e-01 lpdiblc1 = 1.016714599e-07 ppdiblc1 = 5.551115123e-29
+ pdiblc2 = -1.041058628e-02 lpdiblc2 = 2.937964019e-09 ppdiblc2 = -8.673617380e-31
+ pdiblcb = -4.964630236e-01 lpdiblcb = 6.138756232e-8
+ drout = 2.107836980e+00 ldrout = -2.505218234e-7
+ pscbe1 = 8.191380802e+08 lpscbe1 = -4.327808912e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.059378171e-05 lalpha0 = -1.649386622e-12
+ alpha1 = 0.85
+ beta0 = 2.830344734e+01 lbeta0 = -2.075125096e-06 wbeta0 = 5.030914472e-06 pbeta0 = -1.137670875e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.923387179e-01 lkt1 = -1.220746851e-08 wkt1 = -1.289978070e-07 pkt1 = 2.917104808e-14
+ kt2 = 9.136848570e-03 lkt2 = -5.935633008e-9
+ at = -1.610402072e+05 lat = 4.154855845e-02 wat = 1.934967105e-01 pat = -4.375657212e-8
+ ute = 2.035842074e+00 lute = -5.238183671e-7
+ ua1 = 7.768720193e-09 lua1 = -1.216700324e-15
+ ub1 = -6.244158411e-18 lub1 = 1.085443667e-24
+ uc1 = -1.643023312e-10 luc1 = 4.863458112e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.336565660e-06 ltvoff = -2.448291784e-10 wtvoff = -4.463324121e-10 ptvoff = 1.009318263e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.35 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 2.0e-06 wmax = 3.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {1.095894562e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -8.348856930e-08 wvth0 = -1.227781289e-06 pvth0 = 1.633271853e-13
+ k1 = 0.90707349
+ k2 = -1.031447479e-01 lk2 = -4.750730347e-09 wk2 = -5.867975870e-08 pk2 = 9.293768265e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587010672e-01 ldsub = -9.587241274e-12 wdsub = -1.486914722e-10 pdsub = 1.875534753e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-5.542487526e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 4.464083477e-08 wvoff = 5.701931180e-07 pvoff = -8.733006153e-14
+ nfactor = -5.542573853e-01 lnfactor = 4.838451664e-07 wnfactor = 5.894605119e-06 pnfactor = -9.465375898e-13
+ eta0 = 6.941575510e-04 leta0 = -2.367699262e-15 weta0 = -3.672137572e-14 peta0 = 4.631887448e-21
+ etab = -6.517384797e-02 wetab = 4.142593021e-8
+ u0 = 4.935277380e-02 lu0 = -3.258691665e-09 wu0 = -4.056208662e-08 pu0 = 6.374919847e-15
+ ua = -1.262823224e-09 lua = 1.239684637e-17 wua = 1.501679709e-16 pua = -2.425172742e-23
+ ub = 5.317291396e-18 lub = -4.555065233e-25 wub = -6.449707982e-24 pub = 8.910992123e-31
+ uc = 1.532944232e-11 wuc = 1.312871760e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.733684148e+04 lvsat = 3.070605128e-02 wvsat = 4.865111774e-01 pvsat = -6.006969542e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.045636319e+00 lketa = 1.342155556e-07 wketa = 2.081590312e-06 pketa = -2.625634756e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.645277110e+00 lpclm = -1.858255773e-07 wpclm = -2.918923594e-06 ppclm = 3.635272321e-13
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.986056660e+01 lbeta0 = -7.568874690e-07 wbeta0 = -1.173880043e-05 pbeta0 = 1.480685332e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705235600e-01 wkt1 = 5.783321264e-8
+ kt2 = -0.028878939
+ at = 2.915115102e+05 lat = -2.911105650e-02 wat = -4.514923244e-01 pat = 5.694943583e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.943939661e-05 ltvoff = -2.363817788e-10 wtvoff = -2.761606229e-09 ptvoff = 4.624294189e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.36 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.373820865e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.907963906e-08 wvth0 = -8.881784197e-22
+ k1 = 5.401400138e-01 lk1 = 2.262776067e-7
+ k2 = -3.078837623e-02 lk2 = -7.452268871e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.016619280e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.757973648e-7
+ nfactor = 2.421209016e+00 lnfactor = 1.800668548e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.214097967e-02 lu0 = -1.425456455e-8
+ ua = -7.268974247e-10 lua = 4.418949960e-16
+ ub = 1.600068716e-18 lub = -1.153596196e-24
+ uc = 4.074296558e-11 luc = 6.038593027e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.300928259e+00 la0 = 1.609689837e-6
+ ags = 4.247743102e-01 lags = 3.125943624e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.261963924e-25 lb0 = 5.260708209e-29
+ b1 = 0.0
+ keta = -6.319055684e-03 lketa = 1.320733586e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.522173340e-02 lpclm = 1.659870397e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 3.376258697e-03 lpdiblc2 = -1.825262290e-8
+ pdiblcb = 5.959123923e-01 lpdiblcb = -6.207642177e-05 wpdiblcb = -1.665334537e-22 ppdiblcb = 2.930988785e-26
+ drout = 0.56
+ pscbe1 = 6.698134574e+08 lpscbe1 = 2.471094420e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.264125957e-01 lkt1 = 2.012115416e-7
+ kt2 = -4.662013646e-02 lkt2 = 1.110368417e-7
+ at = 140000.0
+ ute = -1.907022139e+00 lute = 2.331657318e-6
+ ua1 = 2.411764120e-10 lua1 = 1.791931074e-15
+ ub1 = -5.160008166e-19 lub1 = 1.814648506e-24 wub1 = 7.703719778e-40
+ uc1 = 1.749127103e-11 luc1 = -4.642332218e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.024741670e-03 ltvoff = 9.902803267e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.37 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.539839+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.55146741
+ k2 = -0.034518962
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.21546827+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.51135
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0314274
+ ua = -7.0477628e-10
+ ub = 1.54232e-18
+ uc = 7.0972e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3815089
+ ags = 0.4404227
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.1073e-24
+ b1 = 0.0
+ keta = -0.0056579
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0024625373
+ pdiblcb = -2.5116166
+ drout = 0.56
+ pscbe1 = 793515780.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.31634
+ kt2 = -0.041061662
+ at = 140000.0
+ ute = -1.7903
+ ua1 = 3.3088e-10
+ ub1 = -4.2516e-19
+ uc1 = 1.5167332e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -0.00052901
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.38 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.287853419e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 8.816548014e-8
+ k1 = 5.483309743e-01 lk1 = 2.501663785e-8
+ k2 = -2.963483658e-02 lk2 = -3.895644861e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.288380869e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.066394782e-7
+ nfactor = 2.558497033e+00 lnfactor = -3.760511442e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.147521304e-02 lu0 = -3.813632729e-10
+ ua = -7.496494897e-10 lua = 3.579148231e-16
+ ub = 1.611793036e-18 lub = -5.541263855e-25
+ uc = 8.123639508e-11 luc = -8.187021115e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.542234158e+00 la0 = -1.281966517e-6
+ ags = 4.269830621e-01 lags = 1.071963796e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.202027848e-24 lb0 = -1.670783420e-29
+ b1 = 0.0
+ keta = -1.059979967e-02 lketa = 3.941726389e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.193698668e-01 lpclm = 3.213592108e-06 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = 1.440006234e-03 lpdiblc2 = 8.155846848e-9
+ pdiblcb = -4.983398045e+00 lpdiblcb = 1.971526497e-5
+ drout = 0.56
+ pscbe1 = 7.870702449e+08 lpscbe1 = 5.141046490e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.141332445e-01 lkt1 = -1.760138183e-8
+ kt2 = -3.996812420e-02 lkt2 = -8.722206193e-9
+ at = 140000.0
+ ute = -1.817437128e+00 lute = 2.164494252e-7
+ ua1 = 3.748619787e-10 lua1 = -3.508062434e-16
+ ub1 = -4.991379884e-19 lub1 = 5.900584965e-25
+ uc1 = 3.254985601e-12 luc1 = 9.501449495e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.840006479e-04 ltvoff = -5.687069897e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.39 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.447262671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.478219384e-8
+ k1 = 5.402698164e-01 lk1 = 5.706889798e-8
+ k2 = -3.270465982e-02 lk2 = -2.675041390e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.136977172e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 4.643930903e-8
+ nfactor = 2.489175018e+00 lnfactor = -1.004173866e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.257575154e-02 lu0 = -4.757254045e-9
+ ua = -5.258090296e-10 lua = -5.321052884e-16
+ ub = 1.379512085e-18 lub = 3.694542658e-25
+ uc = 5.722333245e-11 luc = 1.360899167e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.671868096e-01 la0 = 1.004499947e-6
+ ags = 1.961204884e-01 lags = 1.025137370e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.082155696e-24 lb0 = 8.278934222e-30
+ b1 = 0.0
+ keta = -1.749000880e-03 lketa = 4.225284179e-09 wketa = 1.734723476e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.738214857e-01 lpclm = 5.975541666e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 2.149708243e-03 lpdiblc2 = 5.333975140e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 8.082391335e+08 lpscbe1 = -3.275991519e+1
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.150424779e-01 lkt1 = -1.398614617e-8
+ kt2 = -4.270263241e-02 lkt2 = 2.150570337e-9
+ at = 1.646028932e+05 lat = -9.782444936e-2
+ ute = -1.938283263e+00 lute = 6.969500930e-7
+ ua1 = 2.931550244e-11 lua1 = 1.023133540e-15
+ ub1 = -2.943865257e-19 lub1 = -2.240611654e-25
+ uc1 = 9.646151264e-12 luc1 = 6.960235108e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.929819200e-04 ltvoff = -2.200067937e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.40 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.342389756e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.550650798e-8
+ k1 = 6.302528454e-01 lk1 = -1.207498050e-7
+ k2 = -7.003012197e-02 lk2 = 4.700977557e-08 wk2 = -1.110223025e-22
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.695424173e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.081756878e-8
+ nfactor = 2.927407845e+00 lnfactor = -9.664250529e-7
+ eta0 = 1.556200358e-01 leta0 = -1.494354750e-7
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 3.483318800e-02 lu0 = -9.218255501e-9
+ ua = -1.258399038e-10 lua = -1.322498677e-15
+ ub = 8.990623895e-19 lub = 1.318888206e-24
+ uc = 5.360287210e-11 luc = 2.076351371e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 8.430964044e+04 lvsat = -8.516435621e-3
+ a0 = 1.999457250e+00 la0 = -1.035406831e-6
+ ags = 2.096222212e-01 lags = 9.984561099e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.164311393e-24 lb0 = -4.064934266e-30
+ b1 = 0.0
+ keta = 5.085943942e-02 lketa = -9.973614859e-08 wketa = -2.775557562e-23 pketa = 3.122502257e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.280914582e-01 lpclm = 7.429649702e-7
+ pdiblc1 = 1.649323322e-01 lpdiblc1 = 4.447643207e-7
+ pdiblc2 = 6.380373791e-03 lpdiblc2 = -3.026395354e-09 wpdiblc2 = 1.387778781e-23
+ pdiblcb = -4.921630060e-02 lpdiblcb = 4.785470340e-8
+ drout = 8.528408000e-01 ldrout = -5.786932471e-7
+ pscbe1 = 1.154740475e+09 lpscbe1 = -7.174936905e+02 wpscbe1 = -1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.887283200e-09 lalpha0 = 5.555455173e-14
+ alpha1 = 6.342739440e-01 lalpha1 = 4.263040254e-7
+ beta0 = 1.320696502e+01 lbeta0 = 1.290485941e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.876870551e-01 lkt1 = 1.295694180e-7
+ kt2 = -4.725934087e-02 lkt2 = 1.115524596e-8
+ at = 1.633894479e+05 lat = -9.542651645e-2
+ ute = -1.987865646e+00 lute = 7.949316238e-7
+ ua1 = -5.141762198e-10 lua1 = 2.097147098e-15 pua1 = 1.654361225e-36
+ ub1 = 6.086990610e-19 lub1 = -2.008681104e-24
+ uc1 = 1.034951732e-10 luc1 = -1.158560798e-16 wuc1 = 1.033975766e-31 puc1 = 1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.986982774e-03 ltvoff = 3.570537335e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.41 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.758609527e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.877797783e-9
+ k1 = 4.392858589e-01 lk1 = 6.565994532e-8
+ k2 = -9.358647387e-04 lk2 = -2.043561631e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.934635650e-01 ldsub = 6.494860950e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.017781756e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.351084606e-9
+ nfactor = 1.465327635e+00 lnfactor = 4.607640755e-7
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = -7.632783294e-23 peta0 = 2.879640970e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.774140568e-02 lu0 = -2.295711474e-9
+ ua = -1.371839134e-09 lua = -1.062339720e-16
+ ub = 2.298097091e-18 lub = -4.675993133e-26
+ uc = 7.398743477e-11 luc = 8.654082393e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.364284762e+04 lvsat = 5.070260485e-2
+ a0 = 4.042627414e-01 la0 = 5.217199554e-7
+ ags = 1.278280856e+00 lags = -4.470005522e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.631044528e-02 lketa = 1.463759397e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.355090508e+00 lpclm = -4.547529740e-7
+ pdiblc1 = 7.353854155e-01 lpdiblc1 = -1.120754702e-7
+ pdiblc2 = 5.362028211e-03 lpdiblc2 = -2.032351573e-9
+ pdiblcb = 2.343260119e-02 lpdiblcb = -2.306050500e-08 wpdiblcb = 1.387778781e-23 ppdiblcb = 7.806255642e-30
+ drout = -4.446812800e-01 ldrout = 6.878647659e-07 pdrout = 4.440892099e-28
+ pscbe1 = 5.756251585e+07 lpscbe1 = 3.535012140e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.970567686e-06 lalpha0 = 2.957074856e-12 walpha0 = -1.058791184e-27 palpha0 = 7.411538288e-34
+ alpha1 = 1.281452112e+00 lalpha1 = -2.054298828e-7
+ beta0 = 1.120652299e+01 lbeta0 = 3.243189417e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.318729451e-01 lkt1 = -2.252634408e-8
+ kt2 = -3.479216166e-02 lkt2 = -1.014416479e-9
+ at = 8.375791069e+04 lat = -1.769530623e-2
+ ute = -1.097743715e+00 lute = -7.394843689e-8
+ ua1 = 2.198525948e-09 lua1 = -5.508191447e-16
+ ub1 = -2.277567454e-18 lub1 = 8.087075466e-25
+ uc1 = -7.921055025e-11 luc1 = 6.248955431e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.572253219e-03 ltvoff = -4.777871482e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.42 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.195681646e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.593277925e-8
+ k1 = 3.947279698e-01 lk1 = 8.687556041e-8
+ k2 = 2.918004145e-03 lk2 = -2.227058202e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.095184973e-01 ldsub = 1.049178783e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.946591176e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.274072440e-8
+ nfactor = 2.340878188e+00 lnfactor = 4.388293722e-8
+ eta0 = 0.49
+ etab = -0.000625
+ u0 = 2.832140781e-02 lu0 = -2.571871370e-9
+ ua = -1.145591476e-09 lua = -2.139586271e-16
+ ub = 1.978807687e-18 lub = 1.052652480e-25
+ uc = 7.706502979e-11 luc = -5.999455450e-19
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.071740778e+05 lvsat = 1.093037903e-2
+ a0 = 1.5
+ ags = 2.238075265e+00 lags = -5.016927259e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.163195547e-02 lketa = -1.874083449e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.711604765e-01 lpclm = -3.388206463e-8
+ pdiblc1 = 8.117032664e-01 lpdiblc1 = -1.484131464e-7
+ pdiblc2 = -2.522103509e-04 lpdiblc2 = 6.407895190e-10
+ pdiblcb = 1.559088000e-01 lpdiblcb = -8.613719240e-08 wpdiblcb = 5.551115123e-23 ppdiblcb = 4.163336342e-29
+ drout = 1.0
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.185727360e-06 lalpha0 = 2.584115772e-14
+ alpha1 = 0.85
+ beta0 = 1.701486070e+01 lbeta0 = 4.776307318e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.089088954e-01 lkt1 = 1.415324515e-8
+ kt2 = -5.484301818e-02 lkt2 = 8.532518139e-9
+ at = 6.821312074e+04 lat = -1.029387212e-2
+ ute = -2.132730218e+00 lute = 4.188458967e-7
+ ua1 = -1.764351194e-10 lua1 = 5.799853180e-16
+ ub1 = 2.034441167e-19 lub1 = -3.725913786e-25 pub1 = 3.851859889e-46
+ uc1 = 5.317860243e-11 luc1 = -5.456872969e-19
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.201396422e-03 ltvoff = 2.517790134e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.43 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {7.474055291e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -4.484140953e-08 wvth0 = -3.523114620e-08 pvth0 = 7.967030478e-15
+ k1 = 4.930134021e-01 lk1 = 6.464968589e-8
+ k2 = 3.582618336e-03 lk2 = -2.242087522e-08 wk2 = -3.000113945e-08 pk2 = 6.784337670e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.296581543e-01 ldsub = -5.793162321e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 1.286776183e-02 lcdscd = -1.688729789e-9
+ cit = 0.0
+ voff = {-3.054847668e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.232094461e-08 wvoff = 1.579935062e-07 pvoff = -3.572801952e-14
+ nfactor = 3.337395175e+00 lnfactor = -1.814654281e-07 wnfactor = -1.238110388e-06 pnfactor = 2.799813307e-13
+ eta0 = 1.581403714e+00 leta0 = -2.468056702e-7
+ etab = 9.611909611e-02 letab = -2.187732292e-08 wetab = 4.163336342e-23 petab = -1.301042607e-29
+ u0 = -1.959584230e-02 lu0 = 8.263943902e-09 wu0 = 2.056749245e-08 pu0 = -4.651050472e-15
+ ua = -4.068051533e-09 lua = 4.469148005e-16 wua = -8.573060992e-17 pua = 1.938677720e-23
+ ub = 2.368417726e-18 lub = 1.716039230e-26 wub = 1.998290978e-24 pub = -4.518855286e-31
+ uc = -1.503555767e-10 luc = 5.082804073e-17 wuc = 4.046784666e-16 puc = -9.151236971e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.944225614e+05 lvsat = -8.799644062e-03 wvsat = -1.452665614e-01 pvsat = 3.284999913e-8
+ a0 = 1.5
+ ags = -2.725047683e+00 lags = 6.206480450e-07 wags = 1.554312234e-21 pags = 1.526556659e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.801076620e-01 lketa = 7.692881892e-08 wketa = 4.109482272e-07 pketa = -9.293018831e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.565153056e-01 lpclm = -5.318386426e-08 wpclm = 2.735489883e-07 ppclm = -6.185927401e-14
+ pdiblc1 = -2.942002886e-01 lpdiblc1 = 1.016714599e-7
+ pdiblc2 = -1.041058628e-02 lpdiblc2 = 2.937964019e-9
+ pdiblcb = -4.964630236e-01 lpdiblcb = 6.138756232e-8
+ drout = 2.107836980e+00 ldrout = -2.505218234e-7
+ pscbe1 = 8.191380802e+08 lpscbe1 = -4.327808912e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.059378171e-05 lalpha0 = -1.649386622e-12
+ alpha1 = 0.85
+ beta0 = 3.041889995e+01 lbeta0 = -2.553505086e-06 wbeta0 = 8.924926207e-07 pbeta0 = -2.018247113e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.016961167e-02 lkt1 = -4.887974151e-08 wkt1 = -4.462463104e-07 pkt1 = 1.009123556e-13
+ kt2 = 9.136848570e-03 lkt2 = -5.935633008e-9
+ at = -6.212976870e+04 lat = 1.918134752e-2
+ ute = 2.035842074e+00 lute = -5.238183671e-07 wute = 1.776356839e-21 pute = 2.220446049e-28
+ ua1 = 7.768720193e-09 lua1 = -1.216700324e-15
+ ub1 = -6.244158411e-18 lub1 = 1.085443667e-24
+ uc1 = -1.643023312e-10 luc1 = 4.863458112e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.458720351e-03 ltvoff = -1.254313153e-09 wtvoff = -9.179286604e-09 ptvoff = 2.075767156e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.44 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.68e-06 wmax = 2.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.602109710e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} wvth0 = 1.579507759e-8
+ k1 = 0.90707349
+ k2 = -1.400157524e-01 wk2 = 1.345032383e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-2.265731474e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} wvoff = -7.083277036e-8
+ nfactor = 2.175168474e+00 wnfactor = 5.550784391e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 3.333201484e-02 wu0 = -9.220964231e-9
+ ua = -1.205708445e-09 wua = 3.843535568e-17
+ ub = 2.478324425e-18 wub = -8.958879980e-25
+ uc = 1.751813957e-10 wuc = -1.814283231e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.380637200e+05 wvsat = 6.512693613e-2
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.125962559e-01 wketa = -1.842392267e-7
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.158900541e-01 wpclm = -1.226394245e-7
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.406453525e+01 wbeta0 = -4.001286279e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.432283650e-01 wkt1 = 2.000643140e-7
+ kt2 = -0.028878939
+ at = 60720.487
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.574745046e-03 wtvoff = 4.115322938e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.45 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.333311361e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.151219429e-07 wvth0 = 6.628497158e-09 pvth0 = 2.686800928e-13
+ k1 = 4.509691655e-01 lk1 = 6.516985304e-06 wk1 = 1.459086540e-07 pk1 = -1.029337177e-11
+ k2 = 2.183126725e-03 lk2 = -2.506611043e-06 wk2 = -5.395067680e-08 pk2 = 3.979582397e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.779855702e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 5.556852364e-07 wvoff = -3.874119821e-08 pvoff = -1.360540014e-12
+ nfactor = 2.235792097e+00 lnfactor = -5.452748910e-07 wnfactor = 3.033943685e-07 pnfactor = 3.838625022e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.250559414e-02 lu0 = 1.146096629e-07 wu0 = -5.966120923e-10 pu0 = -2.108582158e-13
+ ua = -7.599440421e-10 lua = -1.379098595e-15 wua = 5.407358511e-17 pua = 2.979659036e-21
+ ub = 1.640904249e-18 lub = 8.142629409e-24 wub = -6.681844800e-26 pub = -1.521124663e-29
+ uc = -7.946279064e-11 luc = 5.618322440e-15 wuc = 1.966905152e-16 puc = -8.205075772e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.024781168e+00 la0 = 1.054946940e-05 wa0 = 4.518545145e-07 pa0 = -1.462800038e-11
+ ags = 3.255317977e-01 lags = 6.609171617e-06 wags = 1.623887370e-07 pags = -1.030297602e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.676380820e-24 lb0 = 3.572977822e-28 wb0 = 1.497228208e-29 pb0 = -4.985599081e-34
+ b1 = 0.0
+ keta = -5.251190380e-03 lketa = -2.467254744e-07 wketa = -1.747328776e-09 pketa = 4.253233787e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.115884910e-02 lpclm = 6.466704889e-07 wpclm = 3.937366444e-08 ppclm = -7.865336756e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 6.519696279e-03 lpdiblc2 = -1.208370063e-07 wpdiblc2 = -5.143550334e-09 ppdiblc2 = 1.678569801e-13
+ pdiblcb = 9.806954753e+00 lpdiblcb = -2.630310212e-04 wpdiblcb = -1.507186282e-05 ppdiblcb = 3.288183938e-10
+ drout = 0.56
+ pscbe1 = 2.884416584e+08 lpscbe1 = 1.194071452e+04 wpscbe1 = 6.240318100e+02 ppscbe1 = -1.549496892e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.383284327e-01 lkt1 = -9.410351868e-07 wkt1 = 1.949766955e-08 pkt1 = 1.869037761e-12
+ kt2 = -4.794737592e-02 lkt2 = -1.044018015e-06 wkt2 = 2.171738047e-09 pkt2 = 1.889995471e-12
+ at = 140000.0
+ ute = -1.881602031e+00 lute = -2.725108706e-05 wute = -4.159446421e-08 pute = 4.840571214e-11
+ ua1 = 7.209456077e-10 lua1 = -6.695541727e-14 wua1 = -7.850376991e-16 pua1 = 1.124900486e-19
+ ub1 = -1.152844987e-18 lub1 = 4.443852500e-23 wub1 = 1.042056652e-24 pub1 = -6.974468188e-29
+ uc1 = -4.396503424e-12 luc1 = 2.680225168e-15 wuc1 = 3.581457136e-17 puc1 = -4.461565845e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.972241333e-03 ltvoff = -1.021736680e-08 wtvoff = 1.550376644e-09 ptvoff = 3.292227211e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.46 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.275681626e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} wvth0 = 2.007855040e-8
+ k1 = 7.772076985e-01 wk1 = -3.693747708e-7
+ k2 = -1.232971485e-01 wk2 = 1.452661486e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.501681166e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} wvoff = -1.068494657e-7
+ nfactor = 2.208495782e+00 wnfactor = 4.955549055e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.824292306e-02 wu0 = -1.115211771e-8
+ ua = -8.289813472e-10 wua = 2.032345157e-16
+ ub = 2.048522089e-18 wub = -8.282893664e-25
+ uc = 2.017889209e-10 wuc = -2.140533730e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.552884771e+00 wa0 = -2.804192535e-7
+ ags = 6.563851527e-01 wags = -3.533754741e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.209850140e-24 wb0 = -9.985492947e-30
+ b1 = 0.0
+ keta = -1.760220133e-02 wketa = 1.954424527e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 4.706282143e-04 wpdiblc2 = 3.259324983e-9
+ pdiblcb = -3.360307483e+00 wpdiblcb = 1.388697615e-6
+ drout = 0.56
+ pscbe1 = 8.861906187e+08 wpscbe1 = -1.516421704e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.854364012e-01 wkt1 = 1.130611976e-7
+ kt2 = -1.002106372e-01 wkt2 = 9.678440342e-8
+ at = 140000.0
+ ute = -3.245784127e+00 wute = 2.381582478e-6
+ ua1 = -2.630824588e-09 wua1 = 4.846183907e-15
+ ub1 = 1.071735633e-18 wub1 = -2.449343380e-24
+ uc1 = 1.297748482e-10 wuc1 = -1.875302159e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.483719969e-03 wtvoff = 3.198456738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.47 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.085196784e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.519333006e-07 wvth0 = 3.316034048e-08 pvth0 = -1.043421367e-13
+ k1 = 8.131687922e-01 lk1 = -2.868305740e-07 wk1 = -4.333493544e-07 pk1 = 5.102699796e-13
+ k2 = -1.314425024e-01 lk2 = 6.496845011e-08 wk2 = 1.665860510e-07 pk2 = -1.700504411e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.640068340e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.103794920e-07 wvoff = -1.060822123e-07 pvoff = -6.119717226e-15
+ nfactor = 2.314597209e+00 lnfactor = -8.462794098e-07 wnfactor = 3.990888915e-07 pnfactor = 7.694260470e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.678175693e-02 lu0 = 1.165445982e-08 wu0 = -8.683002255e-09 pu0 = -1.969400068e-14
+ ua = -1.111259757e-09 lua = 2.251490986e-15 wua = 5.916963713e-16 pua = -3.098424591e-21
+ ub = 2.340001023e-18 lub = -2.324875619e-24 wub = -1.191553621e-24 pub = 2.897445097e-30
+ uc = 2.405632926e-10 luc = -3.092696615e-16 wuc = -2.607037344e-16 puc = 3.720896274e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.764730513e+00 la0 = -1.689710447e-06 wa0 = -3.640667807e-07 pa0 = 6.671840526e-13
+ ags = 6.019451518e-01 lags = 4.342208517e-07 wags = -2.862873180e-07 pags = -5.351042572e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.637072031e-23 lb0 = -6.509221038e-29 wb0 = -1.991141244e-29 pb0 = 7.917048383e-35
+ b1 = 0.0
+ keta = -4.345760672e-03 lketa = -1.057351736e-07 wketa = -1.023337145e-08 pketa = 2.375103206e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.918176595e-01 lpclm = 2.196218356e-06 wpclm = -2.087113809e-07 ppclm = 1.664710358e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.953831242e-03 lpdiblc2 = 2.731395435e-08 wpdiblc2 = 7.189557173e-09 ppdiblc2 = -3.134806646e-14
+ pdiblcb = -6.675716521e+00 lpdiblcb = 2.644415339e-05 wpdiblcb = 2.769110261e-06 ppdiblcb = -1.101035900e-11
+ drout = 0.56
+ pscbe1 = 8.142000026e+08 lpscbe1 = 5.742069444e+02 wpscbe1 = -4.439193428e+01 ppscbe1 = -8.554424690e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.803797996e-01 lkt1 = -4.033214272e-08 wkt1 = 1.083980456e-07 pkt1 = 3.719393489e-14
+ kt2 = -9.612799359e-02 lkt2 = -3.256372064e-08 wkt2 = 9.189338339e-08 pkt2 = 3.901144094e-14
+ at = 140000.0
+ ute = -2.769448426e+00 lute = -3.799318332e-06 wute = 1.557758950e-06 pute = 6.570928497e-12
+ ua1 = -2.166142124e-09 lua1 = -3.706370531e-15 wua1 = 4.157799275e-15 pua1 = 5.490649443e-21
+ ub1 = 7.656477753e-19 lub1 = 2.441398380e-24 wub1 = -2.069546179e-24 pub1 = -3.029314127e-30
+ uc1 = 1.009927653e-10 luc1 = 2.295698080e-16 wuc1 = -1.599265696e-16 puc1 = -2.201704368e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.470842171e-03 ltvoff = -8.078851070e-09 wtvoff = 2.707789518e-09 ptvoff = 3.913628482e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.48 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.539371677e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.865281367e-08 wvth0 = -1.507163089e-08 pvth0 = 8.743474095e-14
+ k1 = 8.258033443e-01 lk1 = -3.370672714e-07 wk1 = -4.672133721e-07 pk1 = 6.449179195e-13
+ k2 = -1.491428103e-01 lk2 = 1.353472816e-07 wk2 = 1.905256497e-07 pk2 = -2.652375414e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.916146277e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.201518345e-07 wvoff = -3.613416191e-08 pvoff = -2.842426785e-13
+ nfactor = 1.279580357e+00 lnfactor = 3.269088357e-06 wnfactor = 1.979237972e-06 pnfactor = -5.513461597e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.958759303e-02 lu0 = 4.980738802e-10 wu0 = -1.147335002e-08 pu0 = -8.599198488e-15
+ ua = -1.332158241e-09 lua = 3.129813399e-15 wua = 1.319414700e-15 pua = -5.991931634e-21
+ ub = 2.992797430e-18 lub = -4.920482916e-24 wub = -2.639789771e-24 pub = 8.655828991e-30
+ uc = 2.316169767e-10 luc = -2.736978929e-16 wuc = -2.853571810e-16 puc = 4.701150836e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = -1.578126545e-01 la0 = 5.954582653e-06 wa0 = 1.840816373e-06 pa0 = -8.099731231e-12
+ ags = 1.361312378e-01 lags = 2.286360324e-06 wags = 9.815933089e-08 pags = -2.063716418e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.111890208e-24 lb0 = 3.225397868e-29 wb0 = 9.866346046e-30 pb0 = -3.922993370e-35
+ b1 = 0.0
+ keta = -8.830851688e-02 lketa = 2.281121641e-07 wketa = 1.416357780e-07 pketa = -3.663420716e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.704547550e-01 lpclm = -3.945323313e-08 wpclm = 1.691371210e-07 ppclm = 1.623333279e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 4.275440790e-03 lpdiblc2 = -1.430614430e-09 wpdiblc2 = -3.478297903e-09 ppdiblc2 = 1.106877615e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.147432962e+09 lpscbe1 = -7.507726199e+02 wpscbe1 = -5.550167553e+02 ppscbe1 = 1.174871265e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.710108522e-01 lkt1 = -7.758435171e-08 wkt1 = 9.158004335e-08 pkt1 = 1.040645990e-13
+ kt2 = -9.784205172e-02 lkt2 = -2.574839239e-08 wkt2 = 9.022363930e-08 pkt2 = 4.565057053e-14
+ at = 1.534436066e+05 lat = -5.345360828e-02 wat = 1.825973975e-02 pat = -7.260320858e-8
+ ute = -2.510701879e+00 lute = -4.828129792e-06 wute = 9.366382773e-07 pute = 9.040588764e-12
+ ua1 = 2.066007674e-09 lua1 = -2.053397370e-14 wua1 = -3.332602741e-15 pua1 = 3.527350655e-20
+ ub1 = -3.516702540e-18 lub1 = 1.946860563e-23 wub1 = 5.272617693e-24 pub1 = -3.222275622e-29
+ uc1 = 5.638247705e-11 luc1 = 4.069463810e-16 wuc1 = -7.647380863e-17 puc1 = -5.519899639e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.542903231e-03 ltvoff = -3.816190495e-09 wtvoff = 3.026992943e-09 ptvoff = 2.644432251e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.49 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.135899949e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 5.107868690e-08 wvth0 = 3.378755544e-08 pvth0 = -9.117656076e-15
+ k1 = 7.232444938e-01 lk1 = -1.343970348e-07 wk1 = -1.521605605e-07 pk1 = 2.233071647e-14
+ k2 = -1.174196140e-01 lk2 = 7.265793141e-08 wk2 = 7.754257277e-08 pk2 = -4.196761574e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-07 wdsub = 8.881784197e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-5.865689744e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.259072270e-08 wvoff = -1.814399801e-07 pvoff = 2.901379841e-15
+ nfactor = 3.081513941e+00 lnfactor = -2.917774696e-07 wnfactor = -2.521610309e-07 pnfactor = -1.103913697e-12
+ eta0 = 1.556201771e-01 leta0 = -1.494357543e-07 weta0 = -2.312722238e-13 peta0 = 4.570253672e-19
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 5.166343878e-02 lu0 = -2.336543963e-08 wu0 = -2.753903640e-08 pu0 = 2.314878273e-14
+ ua = 2.195974806e-09 lua = -3.842257326e-15 wua = -3.799143616e-15 pua = 4.123035722e-21
+ ub = -1.652587243e-18 lub = 4.259428972e-24 wub = 4.175218364e-24 pub = -4.811553926e-30
+ uc = 9.755077482e-11 luc = -8.764844988e-18 wuc = -7.191116217e-17 puc = 4.831672182e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.250579846e+05 lvsat = -8.904070550e-02 wvsat = -6.667578212e-02 pvsat = 1.317604134e-7
+ a0 = 3.837564157e+00 la0 = -1.940825297e-06 wa0 = -3.007661246e-06 pa0 = 1.481519938e-12
+ ags = -2.127519340e-01 lags = 2.975800920e-06 wags = 6.911232273e-07 pags = -3.235493720e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.622378042e-23 lb0 = -1.583661612e-29 wb0 = -1.973269209e-29 pb0 = 1.926179113e-35
+ b1 = 0.0
+ keta = 2.757168205e-01 lketa = -4.912514101e-07 wketa = -3.679300853e-07 pketa = 6.406293751e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.433166066e-01 lpclm = 2.161510450e-06 wpclm = 1.425869331e-06 ppclm = -2.321140435e-12
+ pdiblc1 = -6.318451294e-01 lpdiblc1 = 2.019304947e-06 wpdiblc1 = 1.303752619e-06 ppdiblc1 = -2.576392485e-12
+ pdiblc2 = 1.095896664e-02 lpdiblc2 = -1.463817048e-08 wpdiblc2 = -7.491869069e-09 ppdiblc2 = 1.900013862e-14
+ pdiblcb = -1.882408497e-01 lpdiblcb = 3.225861198e-07 wpdiblcb = 2.274833673e-07 ppdiblcb = -4.495380715e-13
+ drout = 1.240960114e+00 ldrout = -1.345669796e-06 wdrout = -6.350726477e-07 pdrout = 1.254989922e-12
+ pscbe1 = 2.182036796e+09 lpscbe1 = -2.795290502e+03 wpscbe1 = -1.680946478e+03 ppscbe1 = 3.399861523e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -8.291676297e-08 lalpha0 = 2.231388803e-13 walpha0 = 1.387633343e-13 palpha0 = -2.742152203e-19
+ alpha1 = -4.229498316e-01 lalpha1 = 2.515521988e-06 walpha1 = 1.729916234e-06 palpha1 = -3.418549747e-12
+ beta0 = 1.131583479e+01 lbeta0 = 5.027616468e-06 wbeta0 = 3.094422354e-06 pbeta0 = -6.114999413e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.666636745e-01 lkt1 = 3.090522339e-07 wkt1 = 2.928562207e-07 pkt1 = -2.936845010e-13
+ kt2 = -1.852391368e-01 lkt2 = 1.469601338e-07 wkt2 = 2.257738565e-07 pkt2 = -2.222150934e-13
+ at = 2.424843300e+05 lat = -2.294101872e-01 wat = -1.294215318e-01 pat = 2.192350687e-7
+ ute = -8.285966809e+00 lute = 6.584579146e-06 wute = 1.030546957e-05 pute = -9.473496027e-12
+ ua1 = -1.914313411e-08 lua1 = 2.137817490e-14 wua1 = 3.048222847e-14 pua1 = -3.154919874e-20
+ ub1 = 1.585972640e-17 lub1 = -1.882185315e-23 wub1 = -2.495498152e-23 pub1 = 2.751109078e-29
+ uc1 = 6.271597049e-10 luc1 = -7.209870469e-16 wuc1 = -8.568628472e-16 puc1 = 9.901649091e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.039319248e-03 ltvoff = 3.093203066e-09 wtvoff = 6.630765231e-09 ptvoff = -4.477111902e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.50 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.574998711e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 8.216676046e-09 wvth0 = 3.004390735e-08 pvth0 = -5.463346403e-15
+ k1 = 5.557583055e-01 lk1 = 2.909226309e-08 wk1 = -1.905817679e-07 pk1 = 5.983504023e-14
+ k2 = -2.812430428e-02 lk2 = -1.450643502e-08 wk2 = 4.448795424e-08 pk2 = -9.701812613e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.479196217e-01 ldsub = 1.094056921e-07 wdsub = 7.452273465e-08 pdsub = -7.274432412e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-4.097212509e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.985346565e-08 wvoff = -2.631240459e-07 pvoff = 8.263613706e-14
+ nfactor = 3.086945135e+00 lnfactor = -2.970790533e-07 wnfactor = -2.653423526e-06 pnfactor = 1.240045070e-12
+ eta0 = -4.616718742e-01 leta0 = 4.531252395e-07 weta0 = 4.625444475e-13 peta0 = -2.202340631e-19
+ etab = -1.632660008e-01 letab = 7.700834592e-08 wetab = -1.410113851e-09 petab = 1.376462894e-15
+ u0 = 3.061335739e-02 lu0 = -2.817697384e-09 wu0 = -4.699322888e-09 pu0 = 8.541161482e-16
+ ua = -1.576921233e-09 lua = -1.593976788e-16 wua = 3.355721464e-16 pua = 8.699081638e-23
+ ub = 2.541609194e-18 lub = 1.653228380e-25 wub = -3.984544719e-25 pub = -3.470272179e-31
+ uc = 1.055135756e-10 luc = -1.653762153e-17 wuc = -5.158565684e-17 puc = 2.847626436e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.351428253e+04 lvsat = 9.503147307e-02 wvsat = 1.426136432e-01 pvsat = -7.253452915e-8
+ a0 = 2.181910458e+00 la0 = -3.246821177e-07 wa0 = -2.908732961e-06 pa0 = 1.384952477e-12
+ ags = 4.162394974e+00 lags = -1.294937483e-06 wags = -4.719224018e-06 pags = 2.045740998e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -3.995377377e-01 lketa = 1.678888733e-07 wketa = 5.452538204e-07 pketa = -2.507623099e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.766725258e+00 lpclm = -1.264767775e-06 wpclm = -2.309832532e-06 ppclm = 1.325412638e-12
+ pdiblc1 = 1.342014350e+00 lpdiblc1 = 9.254964994e-08 wpdiblc1 = -9.926160061e-07 ppdiblc1 = -3.348244008e-13
+ pdiblc2 = -7.510332783e-03 lpdiblc2 = 3.390377589e-09 wpdiblc2 = 2.106281259e-08 ppdiblc2 = -8.873114118e-15
+ pdiblcb = 3.014816994e-01 lpdiblcb = -1.554496904e-07 wpdiblcb = -4.549667345e-07 ppdiblcb = 2.166260411e-13
+ drout = -1.220919908e+00 ldrout = 1.057459922e-06 wdrout = 1.270145295e-06 pdrout = -6.047619004e-13
+ pscbe1 = -2.092469265e+09 lpscbe1 = 1.377208746e+03 wpscbe1 = 3.518058303e+03 ppscbe1 = -1.675074208e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.165315590e-05 lalpha0 = 1.151726583e-11 walpha0 = 1.420716281e-11 palpha0 = -1.400688641e-17
+ alpha1 = 3.395899663e+00 lalpha1 = -1.212194482e-06 walpha1 = -3.459832468e-06 palpha1 = 1.647350792e-12
+ beta0 = 3.522293653e+00 lbeta0 = 1.263517254e-05 wbeta0 = 1.257356615e-05 pbeta0 = -1.536793292e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.990952945e-01 lkt1 = -4.974449421e-08 wkt1 = -5.363347965e-08 pkt1 = 4.453656913e-14
+ kt2 = -3.097782830e-02 lkt2 = -3.619882884e-09 wkt2 = -6.241325025e-09 pkt2 = 4.263277779e-15
+ at = -2.004109801e+04 lat = 2.685033402e-02 wat = 1.698444496e-01 pat = -7.288922932e-8
+ ute = -1.739299944e+00 lute = 1.941419392e-07 wute = 1.049766909e-06 pute = -4.386714567e-13
+ ua1 = 4.535025217e-09 lua1 = -1.734928828e-15 wua1 = -3.823171697e-15 pua1 = 1.937537360e-21
+ ub1 = -6.407326370e-18 lub1 = 2.913818675e-24 wub1 = 6.757450178e-24 pub1 = -3.444555447e-30
+ uc1 = -3.025200316e-10 luc1 = 1.865068124e-16 wuc1 = 3.653972848e-16 puc1 = -2.029272071e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.667945057e-03 ltvoff = -1.977166511e-10 wtvoff = 1.792860831e-09 ptvoff = 2.453407463e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.51 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.673190327e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.541419697e-09 wvth0 = 8.549431395e-08 pvth0 = -3.186528120e-14
+ k1 = 8.060266948e-01 lk1 = -9.006952671e-08 wk1 = -6.730007004e-07 pk1 = 2.895320610e-13
+ k2 = -1.440667317e-01 lk2 = 4.069792861e-08 wk2 = 2.405084776e-07 pk2 = -1.030342405e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.002345918e-01 ldsub = 2.275608468e-07 wdsub = 3.432152042e-07 pdsub = -2.006784818e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = -3.370010952e-03 lcdscd = 4.175717935e-09 wcdscd = 1.435021106e-08 pcdscd = -6.832652094e-15
+ cit = 0.0
+ voff = {-1.243755665e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.014208466e-08 wvoff = -1.150037095e-07 pvoff = 1.211071257e-14
+ nfactor = 1.157484251e+00 lnfactor = 6.216067341e-07 wnfactor = 1.936366198e-06 pnfactor = -9.453190498e-13
+ eta0 = -7.917257321e-01 leta0 = 6.102757632e-07 weta0 = 2.097264744e-06 peta0 = -9.985832464e-13
+ etab = -1.159631597e-01 letab = 5.448576041e-08 wetab = 1.887257547e-07 petab = -8.915406901e-14
+ u0 = 5.311302491e-02 lu0 = -1.353059908e-08 wu0 = -4.056607680e-08 pu0 = 1.793156889e-14
+ ua = 6.572337766e-10 lua = -1.223159308e-15 wua = -2.949930510e-15 pua = 1.651336909e-21
+ ub = 1.575914872e-18 lub = 6.251246697e-25 wub = 6.592462614e-25 pub = -8.506366142e-31
+ uc = 1.150341124e-10 luc = -2.107069180e-17 wuc = -6.212812636e-17 puc = 3.349591362e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.384488319e+05 lvsat = -1.130436383e-03 wvsat = -5.117431715e-02 pvsat = 1.973489516e-8
+ a0 = 1.5
+ ags = 5.953233758e+00 lags = -2.147620298e-06 wags = -6.079046970e-06 pags = 2.693201659e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.665092979e-01 lketa = 5.693564410e-08 wketa = 2.206973675e-07 pketa = -9.622929862e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.971661992e-01 lpclm = 1.940612477e-07 wpclm = 1.257199110e-06 ppclm = -3.729795390e-13
+ pdiblc1 = 3.313561455e+00 lpdiblc1 = -8.461749024e-07 wpdiblc1 = -4.093745520e-06 ppdiblc1 = 1.141735002e-12
+ pdiblc2 = 1.218033609e-02 lpdiblc2 = -5.985058727e-09 wpdiblc2 = -2.034315196e-08 ppdiblc2 = 1.084175622e-14
+ pdiblcb = 4.747103024e-01 lpdiblcb = -2.379300645e-07 wpdiblcb = -5.216491600e-07 ppdiblcb = 2.483759444e-13
+ drout = -3.010246809e-01 ldrout = 6.194646874e-07 wdrout = 2.128843267e-06 pdrout = -1.013618918e-12
+ pscbe1 = 7.775245680e+08 lpscbe1 = 1.070136230e+01 wpscbe1 = 3.677614484e+01 ppscbe1 = -1.751044650e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.230242466e-05 lalpha0 = 1.111515241e-13 walpha0 = -1.491748770e-11 palpha0 = -1.395918170e-19
+ alpha1 = 0.85
+ beta0 = 2.735601155e+01 lbeta0 = 1.287081431e-06 wbeta0 = -1.692103899e-05 pbeta0 = -1.324489608e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.413124179e-01 lkt1 = 1.797019807e-08 wkt1 = 5.302130068e-08 pkt1 = -6.245611361e-15
+ kt2 = -8.882559683e-02 lkt2 = 2.392352224e-08 wkt2 = 5.560508177e-08 pkt2 = -2.518402296e-14
+ at = 6.449632294e+04 lat = -1.340097544e-02 wat = 6.081729330e-03 pat = 5.084097239e-9
+ ute = -5.002565161e+00 lute = 1.747899986e-06 wute = 4.695859259e-06 pute = -2.174707284e-12
+ ua1 = -6.781547933e-09 lua1 = 3.653299046e-15 wua1 = 1.080782720e-14 pua1 = -5.028807933e-21
+ ub1 = 6.395571014e-18 lub1 = -3.182101674e-24 wub1 = -1.013206578e-23 pub1 = 4.597151125e-30
+ uc1 = 3.765168716e-10 luc1 = -1.368071026e-16 wuc1 = -5.290725897e-16 puc1 = 2.229621011e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.694857120e-03 ltvoff = 1.719641151e-09 wtvoff = 7.352568858e-09 ptvoff = -2.401836395e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.52 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {8.771035309e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -6.651200760e-08 wvth0 = -2.474536520e-07 pvth0 = 4.342624002e-14
+ k1 = -7.060671499e-01 lk1 = 2.518693270e-07 wk1 = 1.962033924e-06 pk1 = -3.063441287e-13
+ k2 = 4.334038736e-01 lk2 = -8.988896420e-08 wk2 = -7.333099227e-07 pk2 = 1.171811572e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.904090211e+00 ldsub = -2.256891467e-07 wdsub = -1.758073834e-06 pdsub = 2.744986161e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 4.418922952e-02 lcdscd = -6.579138468e-09 wcdscd = -5.125075379e-08 pcdscd = 8.002087694e-15
+ cit = 0.0
+ voff = {-1.024407728e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.510233118e-08 wvoff = -1.742437264e-07 pvoff = 2.550701304e-14
+ nfactor = 7.576155152e+00 lnfactor = -8.298858287e-07 wnfactor = -8.173917041e-06 pnfactor = 1.340979961e-12
+ eta0 = 6.158995614e+00 leta0 = -9.615325591e-07 weta0 = -7.490231230e-06 peta0 = 1.169494743e-12
+ etab = 5.018855292e-01 letab = -8.523207072e-08 wetab = -6.639483107e-07 petab = 1.036662334e-13
+ u0 = -8.842795832e-02 lu0 = 1.847691271e-08 wu0 = 1.331962449e-07 pu0 = -2.136234749e-14
+ ua = -1.269058834e-08 lua = 1.795263794e-15 wua = 1.402317116e-14 pua = -2.186892410e-21
+ ub = 1.059986038e-17 lub = -1.415514271e-24 wub = -1.147067046e-23 pub = 1.892374234e-30
+ uc = 3.517486663e-11 luc = -3.011641408e-18 wuc = 1.010983416e-16 puc = -3.415466940e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.833278643e+04 lvsat = 2.150940567e-02 wvsat = 1.101403278e-01 pvsat = -1.674415339e-8
+ a0 = 1.5
+ ags = -1.423642612e+01 lags = 2.417988629e-06 wags = 1.883586134e-05 pags = -2.940956046e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.754556789e-01 lketa = -4.300854788e-08 wketa = -6.617382673e-07 pketa = 1.033211661e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.497935204e+00 lpclm = -2.118758031e-07 wpclm = -1.266879446e-06 ppclm = 1.978054891e-13
+ pdiblc1 = -2.179936755e+00 lpdiblc1 = 3.961028088e-07 wpdiblc1 = 3.085596637e-06 ppdiblc1 = -4.817727165e-13
+ pdiblc2 = -6.490204233e-02 lpdiblc2 = 1.144604200e-08 wpdiblc2 = 8.916338869e-08 ppdiblc2 = -1.392161486e-14
+ pdiblcb = -1.635039818e+00 lpdiblcb = 2.391603887e-07 wpdiblcb = 1.863032714e-06 ppdiblcb = -2.908864758e-13
+ drout = 6.754353698e+00 ldrout = -9.760103575e-07 wdrout = -7.603011667e-06 pdrout = 1.187103830e-12
+ pscbe1 = 8.994074803e+08 lpscbe1 = -1.686075196e+01 wpscbe1 = -1.313433744e+02 ppscbe1 = 2.050742911e-5
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 4.126412212e-05 lalpha0 = -6.438130891e-12 walpha0 = -5.018532593e-11 palpha0 = 7.835736050e-18
+ alpha1 = 0.85
+ beta0 = 7.612893730e+01 lbeta0 = -9.742232906e-06 wbeta0 = -7.390201872e-05 pbeta0 = 1.156096122e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.530414395e-01 lkt1 = 2.062255210e-08 wkt1 = 8.206304986e-08 pkt1 = -1.281299635e-14
+ kt2 = 1.192271299e-01 lkt2 = -2.312468917e-08 wkt2 = -1.801387456e-07 pkt2 = 2.812614319e-14
+ at = -2.477114787e+05 lat = 5.720044798e-02 wat = 3.036640115e-01 pat = -6.220996973e-8
+ ute = 1.175128629e+01 lute = -2.040748965e-06 wute = -1.589720649e-05 pute = 2.482126233e-12
+ ua1 = 3.033529071e-08 lua1 = -4.740154379e-15 wua1 = -3.692527315e-14 pua1 = 5.765364448e-21
+ ub1 = -2.637626537e-17 lub1 = 4.228790318e-24 wub1 = 3.294180424e-23 pub1 = -5.143401546e-30
+ uc1 = -1.066345080e-09 luc1 = 1.894759278e-16 wuc1 = 1.475996313e-15 puc1 = -2.304561604e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.258868818e-03 ltvoff = -9.835266175e-10 wtvoff = -1.048855514e-08 ptvoff = 1.632684021e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.53 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.26e-06 wmax = 1.68e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.511158817e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} wvth0 = 3.067720844e-8
+ k1 = 0.90707349
+ k2 = -1.423055348e-01 wk2 = 1.719705358e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-2.632129917e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} wvoff = -1.087965254e-8
+ nfactor = 2.261007917e+00 wnfactor = 4.146209049e-7
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 2.991062283e-02 wu0 = -3.622602078e-9
+ ua = -1.192511062e-09 wua = 1.684071653e-17
+ ub = 1.533954559e-18 wub = 6.493674149e-25
+ uc = 1.588628867e-11 wuc = 7.922339325e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.760934930e+05 wvsat = 2.899503220e-3
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 0.0
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.14094
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 1.373312271e+01 wbeta0 = 1.421557388e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 1.186386775e+05 wat = -9.477049255e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.040297406e-03 wtvoff = -3.174811500e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.54 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.842573935e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.800276589e-06 wvth0 = -1.769403931e-07 pvth0 = 3.534585356e-12
+ k1 = 4.949059275e-01 lk1 = -4.272885007e-07 wk1 = 9.246916123e-08 pk1 = -1.847176541e-12
+ k2 = -9.994835634e-03 lk2 = 1.224993099e-07 wk2 = -3.913884038e-08 pk2 = 7.818427984e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.652355717e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -3.425783728e-06 wvoff = -1.743104383e-07 pvoff = 3.482049021e-12
+ nfactor = 2.022745174e+00 lnfactor = 1.184954076e-05 wnfactor = 5.625195056e-07 pnfactor = -1.123696615e-11
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.235139522e-02 lu0 = -6.647557703e-07 wu0 = -3.689752273e-08 pu0 = 7.370699321e-13
+ ua = 8.888569869e-10 lua = -3.097786180e-14 wua = -1.951333428e-15 pua = 3.898010194e-20
+ ub = 1.336014698e-18 lub = 6.293741821e-25 wub = 3.040132251e-25 pub = -6.073009531e-30
+ uc = 1.853722886e-10 luc = -3.187657714e-15 wuc = -1.254236246e-16 puc = 2.505479383e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.483199001e+00 la0 = -3.213535043e-06 wa0 = -1.057108436e-07 pa0 = 2.111694188e-12
+ ags = 8.981978616e-01 lags = -1.063429923e-05 wags = -5.341346886e-07 pags = 1.066994718e-11
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.070357563e-09 lb0 = 6.133388025e-14 wb0 = 3.734420637e-15 pb0 = -7.459929453e-20
+ b1 = -1.370788090e-07 lb1 = 2.738304931e-12 wb1 = 1.667264879e-13 pb1 = -3.330550998e-18
+ keta = -1.179579840e-02 lketa = 2.050039111e-07 wketa = 6.212760153e-09 pketa = -1.241069417e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.899094693e-01 lpclm = -6.120257970e-06 wpclm = -3.726426174e-07 ppclm = 7.443959605e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 9.195559666e-03 lpdiblc2 = -1.207594770e-07 wpdiblc2 = -8.398154805e-09 ppdiblc2 = 1.677626825e-13
+ pdiblcb = -1.401431107e+01 lpdiblcb = 2.356337033e-04 wpdiblcb = 1.390151402e-05 ppdiblcb = -2.776985346e-10
+ drout = 0.56
+ pscbe1 = 3.414639747e+09 lpscbe1 = -5.299920474e+04 wpscbe1 = -3.178306654e+03 ppscbe1 = 6.349028596e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.600064000e-01 lkt1 = 3.346530151e-06 wkt1 = 1.674923910e-07 pkt1 = -3.345850783e-12
+ kt2 = -9.922157029e-02 lkt2 = 1.569822975e-06 wkt2 = 6.453561772e-08 pkt2 = -1.289172276e-12
+ at = -2.087443630e+04 lat = 3.213649618e+00 wat = 1.956686811e-01 pat = -3.908704185e-6
+ ute = -5.017918848e+00 lute = 7.451535901e-05 wute = 3.773051226e-06 pute = -7.537098442e-11
+ ua1 = -3.556212340e-09 lua1 = 9.807907904e-14 wua1 = 4.417192524e-15 pua1 = -8.823843859e-20
+ ub1 = 3.672190917e-19 lub1 = -2.615433720e-23 wub1 = -8.067699250e-25 pub1 = 1.611614574e-29
+ uc1 = -6.067838646e-11 luc1 = 7.245357204e-16 wuc1 = 1.042692126e-16 puc1 = -2.082895972e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.790477595e-03 ltvoff = 9.861134827e-08 wtvoff = 4.978146680e-09 ptvoff = -9.944413511e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.55 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.5440763+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.47351598
+ k2 = -0.0038625531
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.23801737+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61593
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0290739
+ ua = -6.6188645e-10
+ ub = 1.367521e-18
+ uc = 2.5799e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3223303
+ ags = 0.3658477
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.0015333577
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.083531
+ pdiblc1 = 0.39
+ pdiblc2 = 0.0031503727
+ pdiblcb = -2.2185512
+ drout = 0.56
+ pscbe1 = 761513800.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.29248
+ kt2 = -0.020636654
+ at = 140000.0
+ ute = -1.2877
+ ua1 = 1.3536e-9
+ ub1 = -9.4206e-19
+ uc1 = -2.4408323e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00014598
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.56 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.357833725e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.614551719e-8
+ k1 = 4.568785944e-01 lk1 = 1.327020504e-7
+ k2 = 5.520842473e-03 lk2 = -7.484323923e-08 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512252687e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.053479967e-7
+ nfactor = 2.642719216e+00 lnfactor = -2.136744325e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.964278566e-02 lu0 = -4.537509378e-9
+ ua = -6.247801648e-10 lua = -2.959647776e-16
+ ub = 1.360332146e-18 lub = 5.733927629e-26
+ uc = 2.621848235e-11 luc = -3.345848257e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.465402906e+00 la0 = -1.141166562e-6
+ ags = 3.665660884e-01 lags = -5.729963354e-9
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.275941100e-02 lketa = 8.954052784e-08 wketa = -1.734723476e-24 pketa = 1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.634155134e-01 lpclm = 3.564906175e-06 wpclm = 1.110223025e-22 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.957262709e-03 lpdiblc2 = 1.540271552e-9
+ pdiblcb = -4.399015674e+00 lpdiblcb = 1.739168118e-5
+ drout = 0.56
+ pscbe1 = 7.777019419e+08 lpscbe1 = -1.291188214e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912573382e-01 lkt1 = -9.752116958e-9
+ kt2 = -2.057529825e-02 lkt2 = -4.893818432e-10
+ at = 140000.0
+ ute = -1.488693675e+00 lute = 1.603152885e-6
+ ua1 = 1.252307935e-09 lua1 = 8.079192830e-16
+ ub1 = -9.358870489e-19 lub1 = -4.923629781e-26
+ uc1 = -3.049530213e-11 luc1 = 4.855057335e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.554421261e-04 ltvoff = -4.861152804e-09 wtvoff = 2.168404345e-25 ptvoff = -8.673617380e-31
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.57 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.415456081e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.323408505e-8
+ k1 = 4.416709045e-01 lk1 = 1.931698936e-7
+ k2 = 7.503140004e-03 lk2 = -8.272512381e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.213233317e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.354617187e-8
+ nfactor = 2.906865782e+00 lnfactor = -1.263957102e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.015445991e-02 lu0 = -6.571995798e-9
+ ua = -2.473648295e-10 lua = -1.796619479e-15
+ ub = 8.224210119e-19 lub = 2.196147102e-24
+ uc = -2.997348756e-12 luc = 1.128202696e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.355665612e+00 la0 = -7.048361580e-7
+ ags = 2.168356558e-01 lags = 5.896186001e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.814126858e-02 lketa = -7.308613666e-08 wketa = 1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.095155328e-01 lpclm = 9.401361739e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.415661641e-03 lpdiblc2 = 7.669887058e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.911105335e+08 lpscbe1 = 2.151803947e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957157780e-01 lkt1 = 7.975246273e-9
+ kt2 = -2.366218282e-02 lkt2 = 1.178449104e-8
+ at = 1.684563584e+05 lat = -1.131463511e-1
+ ute = -1.740618726e+00 lute = 2.604841151e-6
+ ua1 = -6.739841536e-10 lua1 = 8.467118605e-15
+ ub1 = 8.183264192e-19 lub1 = -7.024227620e-24 pub1 = 3.081487911e-45
+ uc1 = -6.492586981e-12 luc1 = -4.688748644e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.417697940e-05 ltvoff = -1.641997133e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.58 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.413693713e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.358235293e-8
+ k1 = 5.981414663e-01 lk1 = -1.160372166e-7
+ k2 = -5.366583585e-02 lk2 = 3.815309147e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.078328123e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.020527275e-8
+ nfactor = 2.874192752e+00 lnfactor = -1.199390751e-6
+ eta0 = 1.556199869e-01 leta0 = -1.494353785e-7
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 2.902145575e-02 lu0 = -4.333025486e-9
+ ua = -9.275965507e-10 lua = -4.523890865e-16
+ ub = 1.780184404e-18 lub = 3.034763837e-25
+ uc = 3.842701720e-11 luc = 3.096008872e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.023864000e+04 lvsat = 1.928977490e-2
+ a0 = 1.364731996e+00 la0 = -7.227525654e-7
+ ags = 3.554742071e-01 lags = 3.156499677e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.678710971e-02 lketa = 3.545980911e-08 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.290014341e-01 lpclm = 2.531204263e-7
+ pdiblc1 = 4.400712671e-01 lpdiblc1 = -9.894763339e-8
+ pdiblc2 = 4.799318577e-03 lpdiblc2 = 9.833207738e-10
+ pdiblcb = -1.209086295e-03 lpdiblcb = -4.701408105e-8
+ drout = 7.188175127e-01 ldrout = -3.138450042e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.117136320e-08 lalpha0 = -2.314772989e-15
+ alpha1 = 9.993488080e-01 lalpha1 = -2.951335560e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.258838054e-01 lkt1 = 6.759137127e-8
+ kt2 = 3.871048534e-04 lkt2 = -3.574017210e-8
+ at = 1.360768260e+05 lat = -4.915999135e-02 wat = -1.164153218e-16
+ ute = 1.869609889e-01 lute = -1.204318517e-6
+ ua1 = 5.918675958e-09 lua1 = -4.560874379e-15
+ ub1 = -4.657704193e-18 lub1 = 3.797153610e-24
+ uc1 = -7.733386419e-11 luc1 = 9.310451173e-17 wuc1 = -5.169878828e-32 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.876515994e-04 ltvoff = -5.877787311e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.59 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.822013033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.724834185e-9
+ k1 = 3.990662161e-01 lk1 = 7.828730192e-8
+ k2 = 8.452701900e-03 lk2 = -2.248304950e-08 pk2 = -6.938893904e-30
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.091905561e-01 ldsub = 4.959692731e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.573068615e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 8.088127714e-9
+ nfactor = 9.053593462e-01 lnfactor = 7.224584146e-7
+ eta0 = -4.616714939e-01 leta0 = 4.531250584e-07 weta0 = 4.510281038e-23 peta0 = 8.153200337e-29
+ etab = -1.644253650e-01 letab = 7.814004309e-8
+ u0 = 2.674967867e-02 lu0 = -2.115462090e-9
+ ua = -1.301021280e-09 lua = -8.787576494e-17
+ ub = 2.214008792e-18 lub = -1.199952198e-25
+ uc = 6.310099629e-11 luc = 6.874929471e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.373948201e+04 lvsat = 3.539519699e-2
+ a0 = -2.095850677e-01 la0 = 8.139949958e-7
+ ags = 2.823539824e-01 lags = 3.870252515e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.875782245e-02 lketa = -3.828231879e-08 wketa = -1.387778781e-23 pketa = 6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.676323403e-01 lpclm = -1.750429920e-7
+ pdiblc1 = 5.259075539e-01 lpdiblc1 = -1.827355231e-07 wpdiblc1 = -4.440892099e-22
+ pdiblc2 = 9.807043116e-03 lpdiblc2 = -3.904899426e-9
+ pdiblcb = -7.258182741e-02 lpdiblcb = 2.265542098e-8
+ drout = -1.766347053e-01 ldrout = 5.602381421e-07 pdrout = 2.220446049e-28
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.765727360e-08 lalpha0 = 1.115456377e-15
+ alpha1 = 5.513023840e-01 lalpha1 = 1.422206881e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.431915482e-01 lkt1 = -1.312751794e-8
+ kt2 = -3.610930687e-02 lkt2 = -1.147107452e-10
+ at = 1.196012296e+05 lat = -3.307756865e-2
+ ute = -8.762049469e-01 lute = -1.665239728e-7
+ ua1 = 1.391698507e-09 lua1 = -1.419287174e-16
+ ub1 = -8.515011762e-19 lub1 = 8.178182225e-26 wub1 = 7.703719778e-40
+ uc1 = -2.098513587e-12 luc1 = 1.966457754e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.193894770e-03 ltvoff = 3.997052018e-12
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.60 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.376105555e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.265750555e-8
+ k1 = 2.527004922e-01 lk1 = 1.479772922e-7
+ k2 = 5.367398760e-02 lk2 = -4.401453159e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.819493130e-01 ldsub = 6.256746383e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413312e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-2.189290578e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.018492623e-8
+ nfactor = 2.749521458e+00 lnfactor = -1.556135568e-7
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.920295691e-02 letab = -1.881473159e-08 wetab = -9.540979118e-24 petab = -3.144186300e-30
+ u0 = 1.976049909e-02 lu0 = 1.212337914e-9
+ ua = -1.768133457e-09 lua = 1.345331586e-16 wua = -1.654361225e-30
+ ub = 2.117932481e-18 lub = -7.424982916e-26
+ uc = 6.395374912e-11 luc = 6.468903149e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.637444689e+04 lvsat = 1.509515535e-2
+ a0 = 1.5
+ ags = 9.551765888e-01 lags = 6.667018692e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.494316756e-02 lketa = -2.218194427e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.364749379e-01 lpclm = -1.125942310e-7
+ pdiblc1 = -5.222503249e-02 lpdiblc1 = 9.253421406e-8
+ pdiblc2 = -4.545350845e-03 lpdiblc2 = 2.928792025e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = -8.673617380e-31
+ pdiblcb = 4.582196898e-02 lpdiblcb = -3.372088902e-8
+ drout = 1.449262890e+00 ldrout = -2.139102352e-7
+ pscbe1 = 8.077610961e+08 lpscbe1 = -3.695337236e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.759816960e-08 lalpha0 = -3.617762081e-15
+ alpha1 = 0.85
+ beta0 = 1.344390976e+01 lbeta0 = 1.981155425e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.977194842e-01 lkt1 = 1.283519537e-8
+ kt2 = -4.310833573e-02 lkt2 = 3.217778860e-9
+ at = 6.949658549e+04 lat = -9.220943808e-3
+ ute = -1.141734153e+00 lute = -4.009595862e-8
+ ua1 = 2.104407137e-09 lua1 = -4.812749535e-16
+ ub1 = -1.934788051e-18 lub1 = 5.975737015e-25 wub1 = -7.703719778e-40 pub1 = 1.925929944e-46
+ uc1 = -5.847484063e-11 luc1 = 4.650737639e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.497385888e-04 ltvoff = -2.550952953e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.61 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {8.578077171e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -7.245201088e-08 wvth0 = -2.239845009e-07 pvth0 = 5.065095909e-14
+ k1 = 0.90707349
+ k2 = -2.063178989e-01 lk2 = 1.477899366e-08 wk2 = 4.477215426e-08 pk2 = -1.012459588e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586410187e-01 ldsub = -2.491733918e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-3.079508919e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 9.946115252e-09 wvoff = 7.571453232e-08 pvoff = -1.712178148e-14
+ nfactor = -4.719921313e+00 lnfactor = 1.533496354e-06 wnfactor = 6.781579434e-06 pnfactor = -1.533559247e-12
+ eta0 = 6.941427212e-04 leta0 = -6.153674857e-16
+ etab = -0.043998
+ u0 = 1.648969595e-02 lu0 = 1.951984255e-09 wu0 = 5.586790544e-09 pu0 = -1.263374466e-15
+ ua = -1.154436704e-09 lua = -4.245770439e-18 wua = -8.042423965e-18 pua = 1.818681586e-24
+ ub = 6.649713698e-20 lub = 3.896535538e-25 wub = 1.340869643e-24 pub = -3.032188976e-31
+ uc = 3.575855327e-10 luc = -5.993181387e-17 wuc = -2.910439482e-16 puc = 6.581551426e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.345212964e+05 lvsat = 6.468779387e-03 wvsat = -6.852025480e-03 pvsat = 1.549489634e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.885609012e-01 lketa = 1.142920518e-07 wketa = 3.891495467e-07 pketa = -8.800072189e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.637956964e-01 lpclm = -2.831803807e-08 wpclm = 1.125540227e-07 ppclm = -2.545251649e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -6.604864909e-08 lalpha0 = 1.982051491e-14 walpha0 = 8.381682544e-14 palpha0 = -1.895400164e-20
+ alpha1 = 0.85
+ beta0 = 1.725522692e+01 lbeta0 = -6.637604737e-07 wbeta0 = -2.294984506e-06 pbeta0 = 5.189786163e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.496479997e-01 lkt1 = 4.719170217e-08 wkt1 = 1.995638701e-07 pkt1 = -4.512857533e-14
+ kt2 = -0.028878939
+ at = 1.660312896e+05 lat = -3.105091565e-02 wat = -1.995638701e-01 pat = 4.512857533e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -9.455125138e-03 ltvoff = 1.736119597e-09 wtvoff = 7.407810858e-09 ptvoff = -1.675172716e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.62 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 1.0e-06 wmax = 1.26e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {1.033117780e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.535196706e-08 wvth0 = 4.537050793e-07 pvth0 = -5.516078120e-14
+ k1 = 0.90707349
+ k2 = -8.384763239e-02 lk2 = -4.343023875e-09 wk2 = -5.390424094e-08 pk2 = 5.282341765e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45862506
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-2.277643275e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.573894174e-09 wvoff = -5.399522478e-08 pvoff = 3.130581154e-15
+ nfactor = 1.596421357e+01 lnfactor = -1.696041731e-06 wnfactor = -1.625234148e-05 pnfactor = 2.062865028e-12
+ eta0 = 0.00069413878
+ etab = -0.043998
+ u0 = 3.128641951e-02 lu0 = -3.583169751e-10 wu0 = -5.295958813e-09 pu0 = 4.358144871e-16
+ ua = -1.178876828e-09 lua = -4.297872073e-19 wua = 2.576422700e-19 pua = 5.227424441e-25
+ ub = 1.121291289e-18 lub = 2.249622141e-25 wub = 1.151282322e-24 pub = -2.736174917e-31
+ uc = -4.773210041e-10 luc = 7.042715317e-17 wuc = 6.791025457e-16 puc = -8.565927871e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.298015183e+05 lvsat = -8.407893334e-03 wvsat = -6.242460122e-02 pvsat = 1.022636932e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 7.465502318e-01 lketa = -9.416686003e-08 wketa = -9.080156090e-07 pketa = 1.145334569e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.824279268e-01 wpclm = -5.046101855e-8
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.907954345e-07 lalpha0 = -2.028209293e-14 walpha0 = -1.955725927e-13 palpha0 = 2.466874455e-20
+ alpha1 = 0.85
+ beta0 = 9.447267864e+00 lbeta0 = 5.553430207e-07 wbeta0 = 5.354963848e-06 pbeta0 = -6.754537199e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.618855327e-01 lkt1 = -4.829069745e-08 wkt1 = -4.656490302e-07 pkt1 = 5.873510608e-14
+ kt2 = -0.028878939
+ at = -3.421257857e+05 lat = 4.829069745e-02 wat = 4.656490302e-01 pat = -5.873510608e-8
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.409281560e-02 ltvoff = -1.940561677e-09 wtvoff = -1.843788106e-08 ptvoff = 2.360270238e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.63 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.546305151e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 5.354570369e-06 wvth0 = 4.264765746e-08 pvth0 = -4.263748003e-12
+ k1 = 7.090279257e-01 lk1 = -1.409865527e-05 wk1 = -1.122918515e-07 pk1 = 1.122650541e-11
+ k2 = -9.771995430e-02 lk2 = 5.618666771e-06 wk2 = 4.475111155e-08 pk2 = -4.474043214e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.595280204e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.287710665e-06 wvoff = 1.025625579e-08 pvoff = -1.025380823e-12
+ nfactor = 2.606060065e+00 lnfactor = 5.908524370e-07 wnfactor = 4.705974636e-09 pnfactor = -4.704851602e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.848989046e-02 lu0 = 6.335997156e-07 wu0 = 5.046444771e-09 pu0 = -5.045240487e-13
+ ua = -1.638741430e-09 lua = 5.847831441e-14 wua = 4.657634413e-16 pua = -4.656522915e-20
+ ub = 1.938728517e-18 lub = -3.419468956e-23 wub = -2.723511518e-25 pub = 2.722861579e-29
+ uc = 8.247136757e-11 luc = -3.392626948e-15 wuc = -2.702132608e-17 puc = 2.701487771e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.422698813e+00 la0 = -6.008447066e-06 wa0 = -4.785560273e-08 pa0 = 4.784418247e-12
+ ags = 3.135876419e-01 lags = 3.128489051e-06 wags = 2.491754151e-08 pags = -2.491159519e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.664903457e-09 lb0 = -9.966755540e-14 wb0 = -7.938242417e-16 pb0 = 7.936348035e-20
+ b1 = 7.433107653e-08 lb1 = -4.449745512e-12 wb1 = -3.544098020e-14 pb1 = 3.543252256e-18
+ keta = -9.043586181e-03 lketa = 4.495913021e-07 wketa = 3.580869151e-09 pketa = -3.580014612e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -8.260293143e-02 lpclm = 9.945419202e-06 wpclm = 7.921248620e-08 ppclm = -7.919358293e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -2.308113044e-03 lpdiblc2 = 3.267660523e-07 wpdiblc2 = 2.602600341e-09 ppdiblc2 = -2.601979257e-13
+ pdiblcb = 3.248672826e+00 lpdiblcb = -3.272891596e-04 wpdiblcb = -2.606766745e-06 ppdiblcb = 2.606144666e-10
+ drout = 0.56
+ pscbe1 = -5.756973567e+08 lpscbe1 = 8.005062783e+04 wpscbe1 = 6.375808926e+02 ppscbe1 = -6.374287403e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.772763127e-01 lkt1 = -9.101514812e-07 wkt1 = -7.249102343e-09 pkt1 = 7.247372418e-13
+ kt2 = -4.277241768e-02 lkt2 = 1.325132363e-06 wkt2 = 1.055430917e-08 pkt2 = -1.055179049e-12
+ at = 2.272342715e+05 lat = -5.222180630e+00 wat = -4.159321017e-02 pat = 4.158328436e-6
+ ute = -8.582581435e-01 lute = -2.570804922e-05 wute = -2.047574318e-07 pute = 2.047085685e-11
+ ua1 = 7.738659558e-10 lua1 = 3.470512042e-14 wua1 = 2.764165910e-16 pua1 = -2.763506269e-20
+ ub1 = -1.341379391e-20 lub1 = -5.559235088e-23 wub1 = -4.427775479e-25 pub1 = 4.426718835e-29
+ uc1 = 1.207163183e-10 luc1 = -8.687721902e-15 wuc1 = -6.919527847e-17 puc1 = 6.917876571e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.830190993e-04 ltvoff = -3.214923601e-08 wtvoff = -2.560596856e-10 ptvoff = 2.559985795e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.64 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {8.413920671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.371430994e-06 wvth0 = -2.843177164e-07 pvth0 = 2.267756773e-12
+ k1 = -3.093204041e-01 lk1 = 6.244009465e-06 wk1 = 7.486123430e-07 pk1 = -5.971033859e-12
+ k2 = 3.081173269e-01 lk2 = -2.488393952e-06 wk2 = -2.983407436e-07 pk2 = 2.379606346e-12
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.665164544e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.703010270e-07 wvoff = -6.837503858e-08 pvoff = 5.453686067e-13
+ nfactor = 2.648737440e+00 lnfactor = -2.616766024e-07 wnfactor = -3.137316424e-08 pnfactor = 2.502366247e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 6.425490847e-02 lu0 = -2.806085081e-07 wu0 = -3.364296514e-08 pu0 = 2.683408654e-13
+ ua = 2.585157423e-09 lua = -2.589886353e-14 wua = -3.105089609e-15 pua = 2.476661701e-20
+ ub = -5.311598759e-19 lub = 1.514413689e-23 wub = 1.815674345e-24 pub = -1.448206551e-29
+ uc = -1.625786688e-10 luc = 1.502525906e-15 wuc = 1.801421739e-16 puc = -1.436838478e-21
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 9.887076327e-01 la0 = 2.661019767e-06 wa0 = 3.190373515e-07 pa0 = -2.544685305e-12
+ ags = 5.395589519e-01 lags = -1.385544570e-06 wags = -1.661169434e-07 pags = 1.324971332e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.534101459e-09 lb0 = 4.414074587e-14 wb0 = 5.292161611e-15 pb0 = -4.221100075e-20
+ b1 = -2.470748182e-07 lb1 = 1.970702352e-12 wb1 = 2.362732013e-13 pb1 = -1.884547187e-18
+ keta = 2.343047201e-02 lketa = -1.991149009e-07 wketa = -2.387246100e-08 pketa = 1.904099956e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.357564328e-01 lpclm = -4.404625155e-06 wpclm = -5.280832413e-07 ppclm = 4.212063752e-12
+ pdiblc1 = 0.39
+ pdiblc2 = 2.129425593e-02 lpdiblc2 = -1.447180802e-07 wpdiblc2 = -1.735066894e-08 ppdiblc2 = 1.383912952e-13
+ pdiblcb = -2.039148028e+01 lpdiblcb = 1.449497539e-04 wpdiblcb = 1.737844497e-05 ppdiblcb = -1.386128405e-10
+ drout = 0.56
+ pscbe1 = 5.206373459e+09 lpscbe1 = -3.545280514e+04 wpscbe1 = -4.250539284e+03 ppscbe1 = 3.390287940e-2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.430167130e-01 lkt1 = 4.030876957e-07 wkt1 = 4.832734896e-08 pkt1 = -3.854655078e-13
+ kt2 = 5.294212413e-02 lkt2 = -5.868743411e-07 wkt2 = -7.036206111e-08 pkt2 = 5.612173686e-13
+ at = -1.499647466e+05 lat = 2.312798254e+00 wat = 2.772880678e-01 pat = -2.211687340e-6
+ ute = -2.715155024e+00 lute = 1.138557540e-05 wute = 1.365049545e-06 pute = -1.088782082e-11
+ ua1 = 3.280622859e-09 lua1 = -1.537019640e-14 wua1 = -1.842777273e-15 pua1 = 1.469824215e-20
+ ub1 = -4.028858998e-18 lub1 = 2.462072861e-23 wub1 = 2.951850319e-24 pub1 = -2.354435960e-29
+ uc1 = -5.067993504e-10 luc1 = 3.847616440e-15 wuc1 = 4.613018565e-16 puc1 = -3.679406344e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.639125827e-03 ltvoff = 1.423824685e-08 wtvoff = 1.707064570e-09 ptvoff = -1.361577917e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.65 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.357833725e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.614551719e-8
+ k1 = 4.568785944e-01 lk1 = 1.327020504e-7
+ k2 = 5.520842473e-03 lk2 = -7.484323923e-08 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512252687e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.053479967e-7
+ nfactor = 2.642719216e+00 lnfactor = -2.136744325e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.964278566e-02 lu0 = -4.537509378e-9
+ ua = -6.247801648e-10 lua = -2.959647776e-16
+ ub = 1.360332146e-18 lub = 5.733927629e-26
+ uc = 2.621848235e-11 luc = -3.345848257e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.465402906e+00 la0 = -1.141166562e-6
+ ags = 3.665660884e-01 lags = -5.729963354e-9
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.275941100e-02 lketa = 8.954052784e-08 wketa = -3.469446952e-24 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.634155134e-01 lpclm = 3.564906175e-06 wpclm = 1.110223025e-22
+ pdiblc1 = 0.39
+ pdiblc2 = 2.957262709e-03 lpdiblc2 = 1.540271552e-9
+ pdiblcb = -4.399015674e+00 lpdiblcb = 1.739168118e-5
+ drout = 0.56
+ pscbe1 = 7.777019419e+08 lpscbe1 = -1.291188214e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912573382e-01 lkt1 = -9.752116958e-9
+ kt2 = -2.057529825e-02 lkt2 = -4.893818432e-10
+ at = 140000.0
+ ute = -1.488693675e+00 lute = 1.603152885e-6
+ ua1 = 1.252307935e-09 lua1 = 8.079192830e-16
+ ub1 = -9.358870489e-19 lub1 = -4.923629781e-26
+ uc1 = -3.049530213e-11 luc1 = 4.855057335e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.554421261e-04 ltvoff = -4.861152804e-09 wtvoff = -2.168404345e-25 ptvoff = -8.673617380e-31
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.66 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.415456081e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.323408505e-8
+ k1 = 4.416709045e-01 lk1 = 1.931698936e-7
+ k2 = 7.503140004e-03 lk2 = -8.272512381e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.213233317e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.354617187e-8
+ nfactor = 2.906865782e+00 lnfactor = -1.263957102e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.015445991e-02 lu0 = -6.571995798e-9
+ ua = -2.473648295e-10 lua = -1.796619479e-15
+ ub = 8.224210119e-19 lub = 2.196147102e-24
+ uc = -2.997348756e-12 luc = 1.128202696e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.355665612e+00 la0 = -7.048361580e-7
+ ags = 2.168356558e-01 lags = 5.896186001e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.814126858e-02 lketa = -7.308613666e-08 wketa = 1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.095155328e-01 lpclm = 9.401361739e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.415661641e-03 lpdiblc2 = 7.669887058e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.911105335e+08 lpscbe1 = 2.151803947e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957157780e-01 lkt1 = 7.975246273e-9
+ kt2 = -2.366218282e-02 lkt2 = 1.178449104e-8
+ at = 1.684563584e+05 lat = -1.131463511e-1
+ ute = -1.740618726e+00 lute = 2.604841151e-6
+ ua1 = -6.739841536e-10 lua1 = 8.467118605e-15 pua1 = -3.308722450e-36
+ ub1 = 8.183264192e-19 lub1 = -7.024227620e-24 pub1 = -3.081487911e-45
+ uc1 = -6.492586981e-12 luc1 = -4.688748644e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.417697940e-05 ltvoff = -1.641997133e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.67 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.413693713e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.358235293e-8
+ k1 = 5.981414663e-01 lk1 = -1.160372166e-7
+ k2 = -5.366583585e-02 lk2 = 3.815309147e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.078328123e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.020527275e-8
+ nfactor = 2.874192752e+00 lnfactor = -1.199390751e-6
+ eta0 = 1.556199869e-01 leta0 = -1.494353785e-7
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 2.902145575e-02 lu0 = -4.333025486e-9
+ ua = -9.275965507e-10 lua = -4.523890865e-16
+ ub = 1.780184404e-18 lub = 3.034763837e-25
+ uc = 3.842701720e-11 luc = 3.096008872e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.023864000e+04 lvsat = 1.928977490e-2
+ a0 = 1.364731996e+00 la0 = -7.227525654e-7
+ ags = 3.554742071e-01 lags = 3.156499677e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.678710971e-02 lketa = 3.545980911e-08 wketa = 1.387778781e-23 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.290014341e-01 lpclm = 2.531204263e-7
+ pdiblc1 = 4.400712671e-01 lpdiblc1 = -9.894763339e-8
+ pdiblc2 = 4.799318577e-03 lpdiblc2 = 9.833207738e-10
+ pdiblcb = -1.209086295e-03 lpdiblcb = -4.701408105e-8
+ drout = 7.188175127e-01 ldrout = -3.138450042e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.117136320e-08 lalpha0 = -2.314772989e-15
+ alpha1 = 9.993488080e-01 lalpha1 = -2.951335560e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.258838054e-01 lkt1 = 6.759137127e-8
+ kt2 = 3.871048534e-04 lkt2 = -3.574017210e-8
+ at = 1.360768260e+05 lat = -4.915999135e-02 wat = -1.164153218e-16
+ ute = 1.869609889e-01 lute = -1.204318517e-6
+ ua1 = 5.918675958e-09 lua1 = -4.560874379e-15
+ ub1 = -4.657704193e-18 lub1 = 3.797153610e-24
+ uc1 = -7.733386419e-11 luc1 = 9.310451173e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.876515994e-04 ltvoff = -5.877787311e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.68 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.822013033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.724834185e-9
+ k1 = 3.990662161e-01 lk1 = 7.828730192e-8
+ k2 = 8.452701900e-03 lk2 = -2.248304950e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.091905561e-01 ldsub = 4.959692731e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.573068615e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 8.088127714e-9
+ nfactor = 9.053593462e-01 lnfactor = 7.224584146e-7
+ eta0 = -4.616714939e-01 leta0 = 4.531250584e-07 weta0 = 5.898059818e-23 peta0 = -1.162264729e-28
+ etab = -1.644253650e-01 letab = 7.814004309e-8
+ u0 = 2.674967867e-02 lu0 = -2.115462090e-9
+ ua = -1.301021280e-09 lua = -8.787576494e-17
+ ub = 2.214008792e-18 lub = -1.199952198e-25
+ uc = 6.310099629e-11 luc = 6.874929471e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.373948201e+04 lvsat = 3.539519699e-2
+ a0 = -2.095850677e-01 la0 = 8.139949958e-7
+ ags = 2.823539824e-01 lags = 3.870252515e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.875782245e-02 lketa = -3.828231879e-08 wketa = -1.387778781e-23 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.676323403e-01 lpclm = -1.750429920e-07 wpclm = 8.881784197e-22
+ pdiblc1 = 5.259075539e-01 lpdiblc1 = -1.827355231e-7
+ pdiblc2 = 9.807043116e-03 lpdiblc2 = -3.904899426e-9
+ pdiblcb = -7.258182741e-02 lpdiblcb = 2.265542098e-8
+ drout = -1.766347053e-01 ldrout = 5.602381421e-07 pdrout = -2.220446049e-28
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.765727360e-08 lalpha0 = 1.115456377e-15
+ alpha1 = 5.513023840e-01 lalpha1 = 1.422206881e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.431915482e-01 lkt1 = -1.312751794e-8
+ kt2 = -3.610930687e-02 lkt2 = -1.147107452e-10
+ at = 1.196012296e+05 lat = -3.307756865e-2
+ ute = -8.762049469e-01 lute = -1.665239728e-7
+ ua1 = 1.391698507e-09 lua1 = -1.419287174e-16
+ ub1 = -8.515011762e-19 lub1 = 8.178182225e-26
+ uc1 = -2.098513587e-12 luc1 = 1.966457754e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.193894770e-03 ltvoff = 3.997052018e-12
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.69 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.376105555e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.265750555e-8
+ k1 = 2.527004922e-01 lk1 = 1.479772922e-7
+ k2 = 5.367398760e-02 lk2 = -4.401453159e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.819493130e-01 ldsub = 6.256746383e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413312e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-2.189290578e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.018492623e-8
+ nfactor = 2.749521458e+00 lnfactor = -1.556135568e-7
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.920295691e-02 letab = -1.881473159e-08 wetab = 1.387778781e-23 petab = 5.854691731e-30
+ u0 = 1.976049909e-02 lu0 = 1.212337914e-9
+ ua = -1.768133457e-09 lua = 1.345331586e-16
+ ub = 2.117932481e-18 lub = -7.424982916e-26
+ uc = 6.395374912e-11 luc = 6.468903149e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.637444689e+04 lvsat = 1.509515535e-2
+ a0 = 1.5
+ ags = 9.551765888e-01 lags = 6.667018692e-8
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 1.494316756e-02 lketa = -2.218194427e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 7.364749379e-01 lpclm = -1.125942310e-7
+ pdiblc1 = -5.222503249e-02 lpdiblc1 = 9.253421406e-8
+ pdiblc2 = -4.545350845e-03 lpdiblc2 = 2.928792025e-09 ppdiblc2 = 4.336808690e-31
+ pdiblcb = 4.582196898e-02 lpdiblcb = -3.372088902e-08 ppdiblcb = -6.938893904e-30
+ drout = 1.449262890e+00 ldrout = -2.139102352e-7
+ pscbe1 = 8.077610961e+08 lpscbe1 = -3.695337236e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.759816960e-08 lalpha0 = -3.617762081e-15
+ alpha1 = 0.85
+ beta0 = 1.344390976e+01 lbeta0 = 1.981155425e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.977194842e-01 lkt1 = 1.283519537e-8
+ kt2 = -4.310833573e-02 lkt2 = 3.217778860e-9
+ at = 6.949658549e+04 lat = -9.220943808e-3
+ ute = -1.141734153e+00 lute = -4.009595862e-8
+ ua1 = 2.104407137e-09 lua1 = -4.812749535e-16
+ ub1 = -1.934788051e-18 lub1 = 5.975737015e-25 wub1 = -7.703719778e-40 pub1 = 1.925929944e-46
+ uc1 = -5.847484063e-11 luc1 = 4.650737639e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.497385888e-04 ltvoff = -2.550952953e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.70 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.235833974e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.948546012e-8
+ k1 = 0.90707349
+ k2 = -1.594989122e-01 lk2 = 4.191535277e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586410187e-01 ldsub = -2.491733918e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-2.287749456e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -7.958416550e-9
+ nfactor = 2.371689147e+00 lnfactor = -7.017206936e-8
+ eta0 = 6.941427212e-04 leta0 = -6.153674857e-16
+ etab = -0.043998
+ u0 = 2.233189578e-02 lu0 = 6.308525528e-10
+ ua = -1.162846800e-09 lua = -2.343944841e-18
+ ub = 1.468666835e-18 lub = 7.257250696e-26
+ uc = 5.323603314e-11 luc = 8.892564569e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.273560193e+05 lvsat = 8.089106481e-3
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.816207447e-01 lketa = 2.226823259e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.814953109e-01 lpclm = -5.493415810e-08 wpclm = -4.440892099e-22
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.16e-8
+ alpha1 = 0.85
+ beta0 = 1.485532343e+01 lbeta0 = -1.210558988e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.24096074
+ kt2 = -0.028878939
+ at = -4.265597014e+04 lat = 1.614078651e-2
+ ute = -1.3190432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.708654057e-03 ltvoff = -1.563638693e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.71 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 8.4e-07 wmax = 1.0e-6
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {3.588940700e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.184207270e-08 wvth0 = 2.092963339e-07 pvth0 = -3.267869240e-14
+ k1 = 0.90707349
+ k2 = -6.431235258e-02 lk2 = -1.067051339e-08 wk2 = -7.258547738e-08 pk2 = 1.133320610e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587284293e-01 ldsub = -1.613967235e-11 wdsub = -9.885022130e-11 pdsub = 1.543407815e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {2.221351670e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -7.836171790e-08 wvoff = -4.842260132e-07 pvoff = 7.560511280e-14
+ nfactor = -5.207334629e+00 lnfactor = 1.113186387e-06 wnfactor = 3.993628981e-06 pnfactor = -6.235492546e-13
+ eta0 = -1.383068870e-02 leta0 = 2.267848679e-09 weta0 = 1.388983239e-08 peta0 = -2.168702870e-15
+ etab = -0.043998
+ u0 = 2.491553369e-02 lu0 = 2.274536641e-10 wu0 = 7.964046169e-10 pu0 = -1.243474313e-16
+ ua = -1.268375502e-09 lua = 1.413288451e-17 wua = 8.584361323e-17 pua = -1.340327840e-23
+ ub = 8.366006974e-18 lub = -1.004350593e-24 wub = -5.776708883e-24 pub = 9.019522181e-31
+ uc = 1.487513236e-10 luc = -6.020810825e-18 wuc = 8.040084801e-17 puc = -1.255346681e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.459714032e+05 lvsat = -1.043102509e-02 wvsat = -7.788757113e-02 pvsat = 1.216105381e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -7.679508232e-01 lketa = 1.138154657e-07 wketa = 5.402744889e-07 pketa = -8.435629760e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 9.659855716e-02 lpclm = 5.162081439e-09 wpclm = 3.161606268e-08 ppclm = -4.936405563e-15
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.371808000e-08 lalpha0 = 5.514423739e-15
+ alpha1 = 0.85
+ beta0 = 1.923203543e+01 lbeta0 = -8.044182041e-07 wbeta0 = -4.002033251e-06 pbeta0 = 6.248614637e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -7.435506831e-01 lkt1 = 7.847238336e-08 wkt1 = 4.002033251e-07 pkt1 = -6.248614637e-14
+ kt2 = -0.028878939
+ at = 4.168356834e+05 lat = -5.560240230e-02 wat = -2.601321613e-01 pat = 4.061599514e-8
+ ute = -2.727950088e-01 lute = -1.633570076e-07 wute = -1.000508313e-06 pute = 1.562153659e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.695413081e-02 ltvoff = 3.926091371e-09 wtvoff = 2.081457494e-08 ptvoff = -3.249904473e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.72 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.73 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.843355012e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.765007359e-7
+ k1 = 6.308143008e-01 lk1 = -1.254632799e-6
+ k2 = -6.654986841e-02 lk2 = 5.000025524e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.523843235e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.145927753e-7
+ nfactor = 2.609337875e+00 lnfactor = 5.257968457e-8
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.200484487e-02 lu0 = 5.638374508e-8
+ ua = -1.314327444e-09 lua = 5.203958101e-15
+ ub = 1.749030239e-18 lub = -3.042969578e-24
+ uc = 6.365044836e-11 luc = -3.019082999e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.389366384e+00 la0 = -5.346889202e-7
+ ags = 3.309432311e-01 lags = 2.784027910e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.111988257e-09 lb0 = -8.869369570e-15
+ b1 = 4.964569199e-08 lb1 = -3.959807912e-13
+ keta = -6.549435865e-03 lketa = 4.000892163e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.742977677e-02 lpclm = 8.850382462e-07 ppclm = -2.220446049e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -4.953474300e-04 lpdiblc2 = 2.907875958e-08 ppdiblc2 = 1.387778781e-29
+ pdiblcb = 1.433005225e+00 lpdiblcb = -2.912531065e-05 wpdiblcb = 5.551115123e-23 ppdiblcb = -6.439293543e-27
+ drout = 0.56
+ pscbe1 = -1.316089196e+08 lpscbe1 = 7.123668276e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.823254642e-01 lkt1 = -8.099395856e-8
+ kt2 = -3.542112043e-02 lkt2 = 1.179229150e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.000875981e+00 lute = -2.287747387e-6
+ ua1 = 9.663958972e-10 lua1 = 3.088392584e-15
+ ub1 = -3.218176240e-19 lub1 = -4.947137544e-24
+ uc1 = 7.252035853e-11 luc1 = -7.731163462e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.046681687e-04 ltvoff = -2.860945615e-09 wtvoff = -4.336808690e-25
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.74 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.357833725e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.614551719e-8
+ k1 = 4.568785944e-01 lk1 = 1.327020504e-7
+ k2 = 5.520842473e-03 lk2 = -7.484323923e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512252687e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.053479967e-7
+ nfactor = 2.642719216e+00 lnfactor = -2.136744325e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.964278566e-02 lu0 = -4.537509378e-9
+ ua = -6.247801648e-10 lua = -2.959647776e-16
+ ub = 1.360332146e-18 lub = 5.733927629e-26
+ uc = 2.621848235e-11 luc = -3.345848257e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.465402906e+00 la0 = -1.141166562e-6
+ ags = 3.665660884e-01 lags = -5.729963354e-9
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.275941100e-02 lketa = 8.954052784e-08 wketa = 3.469446952e-24 pketa = -1.387778781e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.634155134e-01 lpclm = 3.564906175e-06 wpclm = 2.220446049e-22 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 2.957262709e-03 lpdiblc2 = 1.540271552e-9
+ pdiblcb = -4.399015674e+00 lpdiblcb = 1.739168118e-5
+ drout = 0.56
+ pscbe1 = 7.777019419e+08 lpscbe1 = -1.291188214e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.912573382e-01 lkt1 = -9.752116958e-9
+ kt2 = -2.057529825e-02 lkt2 = -4.893818432e-10
+ at = 140000.0
+ ute = -1.488693675e+00 lute = 1.603152885e-6
+ ua1 = 1.252307935e-09 lua1 = 8.079192830e-16
+ ub1 = -9.358870489e-19 lub1 = -4.923629781e-26
+ uc1 = -3.049530213e-11 luc1 = 4.855057335e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.554421261e-04 ltvoff = -4.861152804e-09 wtvoff = 2.168404345e-25 ptvoff = 1.734723476e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.75 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.415456081e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.323408505e-8
+ k1 = 4.416709045e-01 lk1 = 1.931698936e-7
+ k2 = 7.503140004e-03 lk2 = -8.272512381e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.213233317e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.354617187e-8
+ nfactor = 2.906865782e+00 lnfactor = -1.263957102e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.015445991e-02 lu0 = -6.571995798e-9
+ ua = -2.473648295e-10 lua = -1.796619479e-15
+ ub = 8.224210119e-19 lub = 2.196147102e-24
+ uc = -2.997348756e-12 luc = 1.128202696e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.355665612e+00 la0 = -7.048361580e-7
+ ags = 2.168356558e-01 lags = 5.896186001e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.814126858e-02 lketa = -7.308613666e-08 wketa = -1.387778781e-23 pketa = -2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.095155328e-01 lpclm = 9.401361739e-8
+ pdiblc1 = 0.39
+ pdiblc2 = 1.415661641e-03 lpdiblc2 = 7.669887058e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.911105335e+08 lpscbe1 = 2.151803947e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.957157780e-01 lkt1 = 7.975246273e-9
+ kt2 = -2.366218282e-02 lkt2 = 1.178449104e-8
+ at = 1.684563584e+05 lat = -1.131463511e-1
+ ute = -1.740618726e+00 lute = 2.604841151e-6
+ ua1 = -6.739841536e-10 lua1 = 8.467118605e-15
+ ub1 = 8.183264192e-19 lub1 = -7.024227620e-24 pub1 = 3.081487911e-45
+ uc1 = -6.492586981e-12 luc1 = -4.688748644e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.417697940e-05 ltvoff = -1.641997133e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.76 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.413693713e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.358235293e-8
+ k1 = 5.981414663e-01 lk1 = -1.160372166e-7
+ k2 = -5.366583585e-02 lk2 = 3.815309147e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.078328123e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.020527275e-8
+ nfactor = 2.874192752e+00 lnfactor = -1.199390751e-6
+ eta0 = 1.556199869e-01 leta0 = -1.494353785e-7
+ etab = -5.596804500e-02 letab = -2.772905143e-8
+ u0 = 2.902145575e-02 lu0 = -4.333025486e-9
+ ua = -9.275965507e-10 lua = -4.523890865e-16
+ ub = 1.780184404e-18 lub = 3.034763837e-25
+ uc = 3.842701720e-11 luc = 3.096008872e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.023864000e+04 lvsat = 1.928977490e-2
+ a0 = 1.364731996e+00 la0 = -7.227525654e-7
+ ags = 3.554742071e-01 lags = 3.156499677e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.678710971e-02 lketa = 3.545980911e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 4.290014341e-01 lpclm = 2.531204263e-7
+ pdiblc1 = 4.400712671e-01 lpdiblc1 = -9.894763339e-8
+ pdiblc2 = 4.799318577e-03 lpdiblc2 = 9.833207738e-10
+ pdiblcb = -1.209086295e-03 lpdiblcb = -4.701408105e-8
+ drout = 7.188175127e-01 ldrout = -3.138450042e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.117136320e-08 lalpha0 = -2.314772989e-15
+ alpha1 = 9.993488080e-01 lalpha1 = -2.951335560e-7
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.258838054e-01 lkt1 = 6.759137127e-8
+ kt2 = 3.871048534e-04 lkt2 = -3.574017210e-8
+ at = 1.360768260e+05 lat = -4.915999135e-2
+ ute = 1.869609889e-01 lute = -1.204318517e-6
+ ua1 = 5.918675958e-09 lua1 = -4.560874379e-15
+ ub1 = -4.657704193e-18 lub1 = 3.797153610e-24
+ uc1 = -7.733386419e-11 luc1 = 9.310451173e-17 puc1 = -5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.876515994e-04 ltvoff = -5.877787311e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.77 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.034367637e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.782233368e-07 wvth0 = 1.423469851e-07 pvth0 = -1.389500166e-13
+ k1 = -1.877614812e-01 lk1 = 6.511109430e-07 wk1 = 4.672803325e-07 pk1 = -4.561291546e-13
+ k2 = 1.810943869e-01 lk2 = -1.910048134e-07 wk2 = -1.374714662e-07 pk2 = 1.341908472e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.889748954e-01 ldsub = 6.933016149e-08 wdsub = 1.609736674e-08 pdsub = -1.571321918e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {3.837524121e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -6.176729074e-07 wvoff = -5.104639605e-07 pvoff = 4.982822486e-13
+ nfactor = 6.988341140e+00 lnfactor = -5.215359102e-06 wnfactor = -4.843768909e-06 pnfactor = 4.728177207e-12
+ eta0 = -4.616714938e-01 leta0 = 4.531250583e-07 weta0 = -1.059644698e-16 peta0 = 1.034357981e-22
+ etab = -1.664973958e-01 letab = 8.016262691e-08 wetab = 1.649920800e-09 petab = -1.610547090e-15
+ u0 = 4.159403876e-02 lu0 = -1.660557637e-08 wu0 = -1.182029674e-08 pu0 = 1.153821718e-14
+ ua = -1.077074867e-09 lua = -3.064779208e-16 wua = -1.783244976e-16 pua = 1.740689618e-22
+ ub = 1.779380939e-18 lub = 3.042606742e-25 wub = 3.460863361e-25 pub = -3.378273318e-31
+ uc = -1.026813584e-10 luc = 1.687010541e-16 wuc = 1.320095050e-16 puc = -1.288592301e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.380582794e+05 lvsat = -4.373658166e-01 wvsat = -3.856543406e-01 pvsat = 3.764510855e-7
+ a0 = -9.747445963e-01 la0 = 1.560894757e-06 wa0 = 6.092827597e-07 pa0 = -5.947428360e-13
+ ags = -5.943352603e+00 lags = 6.464161575e-06 wags = 4.957418091e-06 pags = -4.839114266e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.213199662e-16 lb0 = -1.184247865e-22 wb0 = -9.660490534e-23 pb0 = 9.429952588e-29
+ b1 = -9.314584709e-18 lb1 = 9.092301459e-24 wb1 = 7.417036141e-24 pb1 = -7.240035991e-30
+ keta = 2.114101305e-01 lketa = -1.970530922e-07 wketa = -1.295171052e-07 pketa = 1.264263090e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.481086146e-01 lpclm = 1.368556195e-07 wpclm = 2.544309914e-07 ppclm = -2.483592502e-13
+ pdiblc1 = -1.973953426e-01 lpdiblc1 = 5.233064731e-07 wpdiblc1 = 5.759530771e-07 ppdiblc1 = -5.622085328e-13
+ pdiblc2 = -5.324133019e-04 lpdiblc2 = 6.187816203e-09 wpdiblc2 = 8.233123035e-09 ppdiblc2 = -8.036647787e-15
+ pdiblcb = -5.340990697e-01 lpdiblcb = 4.731590158e-07 wpdiblcb = 3.674978727e-07 ppdiblcb = -3.587279035e-13
+ drout = -1.766353686e-01 ldrout = 5.602387895e-07 wdrout = 5.281445228e-13 pdrout = -5.155408820e-19
+ pscbe1 = -1.607222313e+09 lpscbe1 = 2.349776360e+03 wpscbe1 = 1.916827798e+03 ppscbe1 = -1.871084619e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.568768658e-05 lalpha0 = -2.504656291e-11 walpha0 = -2.043261945e-11 palpha0 = 1.994501542e-17
+ alpha1 = 5.513023840e-01 lalpha1 = 1.422206881e-7
+ beta0 = 4.142961286e+01 lbeta0 = -2.691169162e-05 wbeta0 = -2.195318647e-05 pbeta0 = 2.142929563e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.974760364e-01 lkt1 = 3.986152520e-08 wkt1 = 4.322576081e-08 pkt1 = -4.219422125e-14
+ kt2 = -3.855180350e-02 lkt2 = 2.269498146e-09 wkt2 = 1.944916102e-09 pkt2 = -1.898502624e-15
+ at = -1.421385482e+05 lat = 2.224160511e-01 wat = 2.084186737e-01 pat = -2.034449705e-7
+ ute = -1.435378758e+00 lute = 3.793057145e-07 wute = 4.452600407e-07 pute = -4.346343550e-13
+ ua1 = -3.451243119e-10 lua1 = 1.553446562e-15 wua1 = 1.383000748e-15 pua1 = -1.349996818e-21
+ ub1 = -5.341608751e-19 lub1 = -2.279854699e-25 wub1 = -2.526923696e-25 pub1 = 2.466621189e-31
+ uc1 = -2.239642498e-10 luc1 = 2.362357099e-16 wuc1 = 1.766676922e-16 puc1 = -1.724516944e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.666561234e-03 ltvoff = -7.668877030e-09 wtvoff = -6.259139628e-09 ptvoff = 6.109771520e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.78 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {8.507765988e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -3.477126297e-08 wvth0 = -1.697402833e-07 pvth0 = 9.645966980e-15
+ k1 = 1.426355886e+00 lk1 = -1.174284437e-07 wk1 = -9.345606642e-07 pk1 = 2.113378102e-13
+ k2 = -3.005643829e-01 lk2 = 3.833026666e-08 wk2 = 2.820736381e-07 pk2 = -6.556968064e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.223806346e-01 ldsub = 5.342448646e-08 wdsub = -3.219473359e-08 pdsub = 7.280388301e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413304e-03 lcdscd = -1.441936597e-09 wcdscd = 6.155763399e-18 pcdscd = -2.930981846e-24
+ cit = 0.0
+ voff = {-9.626290449e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.338777399e-08 wvoff = 5.921949131e-07 pvoff = -2.673333688e-14
+ nfactor = -2.027672734e+00 lnfactor = -9.225103195e-07 wnfactor = 3.803993746e-06 pnfactor = 6.106660880e-13
+ eta0 = 9.325986799e-01 leta0 = -2.107371651e-07 weta0 = -5.891998001e-17 peta0 = 8.103628879e-23
+ etab = 4.334701840e-02 letab = -1.975185307e-08 wetab = -3.299841571e-09 petab = 7.462129661e-16
+ u0 = 9.113687381e-03 lu0 = -1.140511790e-09 wu0 = 8.477864525e-09 pu0 = 1.873531868e-15
+ ua = -2.216026280e-09 lua = 2.358178492e-16 wua = 3.566489928e-16 pua = -8.065117599e-23
+ ub = 2.987188189e-18 lub = -2.708198382e-25 wub = -6.921726734e-25 pub = 1.565251600e-31
+ uc = 3.955184586e-10 luc = -6.850981403e-17 wuc = -2.640190100e-16 puc = 5.970420287e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.760245471e+05 lvsat = 1.407027240e-01 wvsat = 6.150474157e-01 pvsat = -1.000190460e-7
+ a0 = 3.030319055e+00 la0 = -3.460602291e-07 wa0 = -1.218565517e-06 pa0 = 2.755615313e-13
+ ags = 1.340658976e+01 lags = -2.749042582e-06 wags = -9.914836182e-06 pags = 2.242101395e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -2.426399324e-16 lb0 = 5.486962376e-23 wb0 = 1.932098107e-22 pb0 = -4.369169375e-29
+ b1 = 1.862916942e-17 lb1 = -4.212725855e-24 wb1 = -1.483407228e-23 pb1 = 3.354517770e-30
+ keta = -3.103614485e-01 lketa = 5.138114037e-08 wketa = 2.590342103e-07 pketa = -5.857696016e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.375522390e+00 lpclm = -2.571058657e-07 wpclm = -5.088619830e-07 ppclm = 1.150720135e-13
+ pdiblc1 = 1.394380761e+00 lpdiblc1 = -2.345954338e-07 wpdiblc1 = -1.151906154e-06 ppdiblc1 = 2.604874502e-13
+ pdiblc2 = 1.613356198e-02 lpdiblc2 = -1.747454603e-09 wpdiblc2 = -1.646624606e-08 ppdiblc2 = 3.723611017e-15
+ pdiblcb = 9.688564536e-01 lpdiblcb = -2.424522152e-07 wpdiblcb = -7.349957455e-07 ppdiblcb = 1.662089979e-13
+ drout = 1.449264214e+00 ldrout = -2.139105341e-07 wdrout = -1.054410701e-12 pdrout = 2.379706321e-19
+ pscbe1 = 5.622205722e+09 lpscbe1 = -1.092414587e+03 wpscbe1 = -3.833655595e+03 ppscbe1 = 8.669275417e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.128246043e-05 lalpha0 = 1.160169501e-11 walpha0 = 4.086523891e-11 palpha0 = -9.241101665e-18
+ alpha1 = 0.85
+ beta0 = -4.169531597e+01 lbeta0 = 1.266707949e-05 wbeta0 = 4.390637294e-05 pbeta0 = -9.928811551e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.891505079e-01 lkt1 = -1.171615863e-08 wkt1 = -8.645152155e-08 pkt1 = 1.954980126e-14
+ kt2 = -3.822334249e-02 lkt2 = 2.113106030e-09 wkt2 = -3.889832193e-09 pkt2 = 8.796310899e-16
+ at = 5.929761411e+05 lat = -1.275985166e-01 wat = -4.168373475e-01 pat = 9.426193042e-8
+ ute = -2.338653081e-02 lute = -2.929946166e-07 wute = -8.905200814e-07 pute = 2.013786492e-13
+ ua1 = 5.578052773e-09 lua1 = -1.266791282e-15 wua1 = -2.766001494e-15 pua1 = 6.254925134e-22
+ ub1 = -2.569468657e-18 lub1 = 7.410978359e-25 wub1 = 5.053847423e-25 pub1 = -1.142856848e-31
+ uc1 = 3.852566319e-10 luc1 = -5.383628390e-17 wuc1 = -3.533353844e-16 puc1 = 7.990185051e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.173751430e-03 ltvoff = -2.031277919e-09 wtvoff = 3.602389993e-09 ptvoff = 1.414342252e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.79 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {9.940916173e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -6.717994799e-08 wvth0 = -2.950290264e-07 pvth0 = 3.797826219e-14
+ k1 = 9.070734930e-01 lk1 = -4.748850202e-16 wk1 = -2.421877809e-15 pk1 = 3.781419622e-22
+ k2 = -2.067272334e-01 lk2 = 1.711030903e-08 wk2 = 3.760706210e-08 pk2 = -1.028698700e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.587177398e-01 ldsub = -1.984115670e-11 wdsub = -6.109158814e-11 pdsub = 1.381503307e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000031e-03 lcdscd = -5.025100128e-18 wcdscd = -2.450002701e-17 pcdscd = 4.001398171e-24
+ cit = 0.0
+ voff = {-1.030135548e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.865342465e-08 wvoff = 6.381090235e-07 pvoff = -3.711617014e-14
+ nfactor = -7.020338813e+00 lnfactor = 2.065112169e-07 wnfactor = 7.478702808e-06 pnfactor = -2.203179205e-13
+ eta0 = -1.008629497e-02 leta0 = 2.437844358e-09 weta0 = 8.584268489e-09 peta0 = -1.941212071e-15
+ etab = -4.399799987e-02 letab = -2.050434822e-17 wetab = -1.045705744e-16 petab = 1.632724511e-23
+ u0 = 2.439907920e-02 lu0 = -4.597089155e-09 wu0 = -1.646060949e-09 pu0 = 4.162915879e-15
+ ua = -1.214258677e-09 lua = 9.282130514e-18 wua = 4.093835200e-17 pua = -9.257634536e-24
+ ub = 2.675122220e-18 lub = -2.002504882e-25 wub = -9.606787065e-25 pub = 2.172440403e-31
+ uc = -4.621647650e-10 luc = 1.254432394e-16 wuc = 4.104043783e-16 puc = -9.280720448e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.768222694e+05 lvsat = 5.042871777e-02 wvsat = 3.218398961e-01 pvsat = -3.371427036e-8
+ a0 = 1.500000009e+00 la0 = -1.450684017e-15 wa0 = -7.398387680e-15 pa0 = 1.155153306e-21
+ ags = 1.250000002e+00 lags = -3.106048752e-16 wags = -1.584059106e-15 pags = 2.473292682e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 4.747288614e-03 lketa = -1.987628900e-08 wketa = -1.484015103e-07 pketa = 3.355892394e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.253453660e+00 lpclm = -2.295017314e-07 wpclm = -6.146965380e-07 ppclm = 1.390050164e-13
+ pdiblc1 = 3.569721484e-01 lpdiblc1 = 2.483540040e-16 wpdiblc1 = 1.266587724e-15 ppdiblc1 = -1.977599196e-22
+ pdiblc2 = 8.406112143e-03 lpdiblc2 = -6.658944229e-18 wpdiblc2 = -3.396011250e-17 ppdiblc2 = 5.302397410e-24
+ pdiblcb = -1.032957699e-01 lpdiblcb = -1.971667274e-17 wpdiblcb = -1.005533434e-16 ppdiblcb = 1.569999686e-23
+ drout = 5.033266684e-01 ldrout = -1.315386911e-15 wdrout = -6.708376077e-15 pdrout = 1.047419040e-21
+ pscbe1 = 7.914198808e+08 lpscbe1 = -1.299495697e-07 wpscbe1 = -6.627311707e-07 ppscbe1 = 1.034765244e-13
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.520576188e-07 lalpha0 = -2.950116442e-14 walpha0 = -1.038810536e-13 palpha0 = 2.349124621e-20
+ alpha1 = 0.85
+ beta0 = 1.148724706e+01 lbeta0 = 6.405874201e-07 wbeta0 = 2.681938591e-06 pbeta0 = -6.064828653e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -9.585292216e-02 lkt1 = -3.281410148e-08 wkt1 = -1.155467434e-07 pkt1 = 2.612927835e-14
+ kt2 = -2.887893895e-02 lkt2 = -7.882083874e-18 wkt2 = -4.019806710e-17 pkt2 = 6.276368314e-24
+ at = -1.513706568e+05 lat = 4.072509088e-02 wat = 8.656754808e-02 pat = -1.957603905e-8
+ ute = -1.268048809e+00 lute = -1.153166767e-08 wute = -4.060591577e-08 pute = 9.182459393e-15
+ ua1 = -2.384732647e-11 lua1 = -1.487216600e-24 wua1 = -7.584694177e-24 pua1 = 1.184243813e-30
+ ub1 = 7.077531835e-19 lub1 = -2.112662719e-33 wub1 = -1.077442402e-32 pub1 = 1.682275540e-39
+ uc1 = 1.471862498e-10 luc1 = 3.058996623e-26 wuc1 = 1.560062635e-25 puc1 = -2.435824599e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.360570470e-02 ltvoff = -1.245097346e-10 wtvoff = 9.473407279e-09 ptvoff = 8.669388703e-17
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.80 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 7.4e-07 wmax = 8.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {9.709350209e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -6.356436965e-08 wvth0 = -2.780608585e-07 pvth0 = 3.532892033e-14
+ k1 = 0.90707349
+ k2 = -3.683712279e-02 lk2 = -9.415653282e-09 wk2 = -9.446350831e-08 pk2 = 1.033398358e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.584252728e-01 ldsub = 2.582347576e-11 wdsub = 1.425478955e-10 pdsub = -1.798042135e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999993e-03 lcdscd = 8.702153581e-19 wcdscd = 5.565652106e-18 pcdscd = -6.929378946e-25
+ cit = 0.0
+ voff = {-3.340319761e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.993563469e-07 wvoff = 2.352492722e-06 pvoff = -3.047931833e-13
+ nfactor = -3.755233940e+01 lnfactor = 4.973655660e-06 wnfactor = 2.974937407e-05 pnfactor = -3.697571449e-12
+ eta0 = 2.876702308e-02 leta0 = -3.628556861e-09 weta0 = -2.002995755e-08 peta0 = 2.526498726e-15
+ etab = -0.043998
+ u0 = -1.245973038e-01 lu0 = 1.866661010e-08 wu0 = 1.198507859e-07 pu0 = -1.480711580e-14
+ ua = -1.029853534e-09 lua = -1.951015083e-17 wua = -1.040871361e-16 pua = 1.338606508e-23
+ ub = -3.284610577e-18 lub = 7.302783517e-25 wub = 3.500468162e-24 pub = -4.793015873e-31
+ uc = 1.452323505e-09 luc = -1.734773010e-16 wuc = -9.576102154e-16 puc = 1.207891221e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.941120380e+05 lvsat = 1.155826731e-01 wvsat = 6.706839516e-01 pvsat = -8.818138581e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.243131449e-01 lketa = 6.272909085e-08 wketa = 3.462701911e-07 pketa = -4.367713683e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.768628110e-01 lpclm = 1.187309611e-07 wpclm = 8.863940278e-07 ppclm = -9.536926020e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.181192019e-07 lalpha0 = 4.391036365e-14 walpha0 = 2.423891341e-13 palpha0 = -3.057399582e-20
+ alpha1 = 0.85
+ beta0 = 1.955789333e+01 lbeta0 = -6.195310072e-07 wbeta0 = -4.261508034e-06 pbeta0 = 4.776391168e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.541912705e-01 lkt1 = 2.313541487e-08 wkt1 = 1.697916332e-07 pkt1 = -1.842231442e-14
+ kt2 = -0.028878939
+ at = 3.438198224e+05 lat = -3.659196977e-02 wat = -2.019909455e-01 pat = 2.547832990e-8
+ ute = -2.275028667e+00 lute = 1.456941394e-07 wute = 5.938343087e-07 pute = -8.987649950e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.652296395e-02 ltvoff = 6.576419456e-09 wtvoff = 4.435970453e-08 ptvoff = -5.360313021e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.81 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.82 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.318345185e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.525267507e-06 wvth0 = 3.655548926e-08 pvth0 = -7.302374251e-13
+ k1 = 7.553195353e-01 lk1 = -3.741766297e-06 wk1 = -8.669075371e-08 pk1 = 1.731746286e-12
+ k2 = -1.258783113e-01 lk2 = 1.685155596e-06 wk2 = 4.130932686e-08 pk2 = -8.252007314e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.404178983e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.244501636e-07 wvoff = -8.332006530e-09 pvoff = 1.664412956e-13
+ nfactor = 2.680934398e+00 lnfactor = -1.377642201e-06 wnfactor = -4.985137040e-08 pnfactor = 9.958377549e-13
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.632503313e-02 lu0 = 1.698444369e-07 wu0 = 3.954750679e-09 pu0 = -7.900063740e-14
+ ua = -1.802840015e-09 lua = 1.496255165e-14 wua = 3.401425097e-16 pua = -6.794733032e-21
+ ub = 2.179925653e-18 lub = -1.165059497e-23 wub = -3.000247207e-25 pub = 5.993334623e-30
+ uc = 6.597431300e-11 luc = -3.483301360e-16 wuc = -1.618065118e-18 puc = 3.232268885e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.378932276e+00 la0 = -3.262557707e-07 wa0 = 7.265081203e-09 pa0 = -1.451282502e-13
+ ags = 3.988336604e-01 lags = -1.077785658e-06 wags = -4.727088389e-08 pags = 9.442896054e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.789356740e-09 lb0 = -2.240057450e-14 wb0 = -4.716394818e-16 pb0 = 9.421534431e-21
+ b1 = 4.059089170e-07 lb1 = -7.512743427e-12 wb1 = -2.480596709e-13 pb1 = 4.955273721e-18
+ keta = -3.274795282e-02 lketa = 5.633540592e-07 wketa = 1.824155578e-08 pketa = -3.643957991e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.467841810e-01 lpclm = 3.269278057e-06 wpclm = 8.310432329e-08 ppclm = -1.660103264e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -7.548456606e-03 lpdiblc2 = 1.699726277e-07 wpdiblc2 = 4.910952963e-09 ppdiblc2 = -9.810186428e-14
+ pdiblcb = 1.125480882e+01 lpdiblcb = -2.253269950e-04 wpdiblcb = -6.838745051e-06 ppdiblcb = 1.366117012e-10
+ drout = 0.56
+ pscbe1 = -5.189850205e+08 lpscbe1 = 1.486194595e+04 wpscbe1 = 2.697230063e+02 ppscbe1 = -5.388023456e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.763255054e-01 lkt1 = -2.008499515e-07 wkt1 = -4.177663310e-09 pkt1 = 8.345357045e-14
+ kt2 = -3.512857767e-02 lkt2 = 1.120790409e-07 wkt2 = -2.036922630e-10 pkt2 = 4.068984347e-15
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -8.996826457e-01 lute = -4.309199207e-06 wute = -7.045909762e-08 pute = 1.407500517e-12
+ ua1 = 5.387868935e-10 lua1 = 1.163036820e-14 wua1 = 2.977364523e-16 pua1 = -5.947623864e-21
+ ub1 = 8.810493406e-20 lub1 = -1.313580631e-23 wub1 = -2.854216986e-25 pub1 = 5.701622668e-30
+ uc1 = 9.414572346e-11 luc1 = -1.205107577e-15 wuc1 = -1.505735234e-17 puc1 = 3.007877181e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 2.617593890e-04 ltvoff = 1.991433202e-09 wtvoff = 1.691330109e-10 ptvoff = -3.378624028e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.83 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.205292633e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.021256004e-08 wvth0 = -5.900703830e-08 pvth0 = 3.198229128e-14
+ k1 = 5.911392919e-01 lk1 = -2.432242347e-06 wk1 = -9.348330698e-08 pk1 = 1.785924615e-12
+ k2 = -3.965644413e-02 lk2 = 9.974382572e-07 wk2 = 3.145613147e-08 pk2 = -7.466103049e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.507799660e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.180090212e-08 wvoff = -3.100562950e-10 pvoff = 1.024571295e-13
+ nfactor = 1.570736561e+00 lnfactor = 7.477446735e-06 wnfactor = 7.464022270e-07 pnfactor = -5.355189229e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 5.414455187e-02 lu0 = -1.318091880e-07 wu0 = -1.706013878e-08 pu0 = 8.861697893e-14
+ ua = 1.746990347e-09 lua = -1.335137810e-14 wua = -1.651421116e-15 pua = 9.090249297e-21
+ ub = -4.422287084e-19 lub = 9.264064832e-24 wub = 1.255090677e-24 pub = -6.410477284e-30
+ uc = 1.381727663e-10 luc = -9.241948184e-16 wuc = -7.795175273e-17 puc = 6.411705627e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.842239813e+00 la0 = -4.021659693e-06 wa0 = -2.623847553e-07 pa0 = 2.005635518e-12
+ ags = 4.042621016e-01 lags = -1.121083643e-06 wags = -2.624705547e-08 pags = 7.766006907e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.158989107e-08 lb0 = -4.993777692e-13 wb0 = -4.288393253e-14 pb0 = 3.477077519e-19
+ b1 = -7.802471032e-07 lb1 = 1.948198308e-12 wb1 = 5.432720135e-13 pb1 = -1.356495415e-18
+ keta = 1.893225442e-02 lketa = 1.511456978e-07 wketa = -2.206633618e-08 pketa = -4.289457096e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.867328499e+00 lpclm = -1.279555860e-05 wpclm = -1.553226902e-06 ppclm = 1.139149713e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 3.394918562e-02 lpdiblc2 = -1.610182104e-07 wpdiblc2 = -2.157911807e-08 ppdiblc2 = 1.131865449e-13
+ pdiblcb = -3.386442646e+01 lpdiblcb = 1.345501618e-04 wpdiblcb = 2.051623515e-05 ppdiblcb = -8.157534117e-11
+ drout = 0.56
+ pscbe1 = 1.711985740e+09 lpscbe1 = -2.932580246e+03 wpscbe1 = -6.505249915e+02 ppscbe1 = 1.951999728e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.248595398e-01 lkt1 = 1.862641072e-07 wkt1 = 2.339660812e-08 pkt1 = -1.364825686e-13
+ kt2 = -9.319538423e-02 lkt2 = 5.752277871e-07 wkt2 = 5.056405871e-08 pkt2 = -4.008615018e-13
+ at = 140000.0
+ ute = -3.224607310e+00 lute = 1.423471610e-05 wute = 1.208685418e-06 pute = -8.795130101e-12
+ ua1 = -5.233895304e-10 lua1 = 2.010243181e-14 wua1 = 1.236386183e-15 pua1 = -1.343442177e-20
+ ub1 = -3.190224405e-19 lub1 = -9.888503004e-24 wub1 = -4.295117233e-25 pub1 = 6.850904301e-30
+ uc1 = 2.437299205e-10 luc1 = -2.398211476e-15 wuc1 = -1.909380865e-16 puc1 = 1.703636373e-21
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.418437929e-04 ltvoff = -1.040171694e-09 wtvoff = 7.909647466e-11 ptvoff = -2.660480370e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.84 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.013446296e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 9.649327279e-08 wvth0 = -4.163698229e-08 pvth0 = -3.708341376e-14
+ k1 = -3.497273802e-01 lk1 = 1.308771499e-06 wk1 = 5.510363804e-07 pk1 = -7.767733172e-13
+ k2 = 3.190818100e-01 lk2 = -4.289538298e-07 wk2 = -2.169466195e-07 pk2 = 2.410728159e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.436826144e+00 ldsub = 7.939652317e-06 wdsub = 1.390354101e-06 pdsub = -5.528236994e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.079761844e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -6.096081592e-07 wvoff = -7.892157842e-08 pvoff = 4.150272327e-13
+ nfactor = 6.511345077e+00 lnfactor = -1.216708465e-05 wnfactor = -2.509734052e-06 pnfactor = 7.591651452e-12
+ eta0 = -4.491589281e-01 leta0 = 2.104007864e-06 weta0 = 3.684438368e-07 peta0 = -1.464982803e-12
+ etab = 3.925980567e-01 letab = -1.839352787e-06 wetab = -3.220987001e-07 petab = 1.280708237e-12
+ u0 = 3.066007229e-02 lu0 = -3.843170330e-08 wu0 = -3.520487959e-10 pu0 = 2.218334086e-14
+ ua = 2.838977358e-09 lua = -1.769326696e-14 wua = -2.148964511e-15 pua = 1.106854950e-20
+ ub = -4.919382610e-18 lub = 2.706583764e-23 wub = 3.997914510e-24 pub = -1.731631787e-29
+ uc = -2.628408164e-10 luc = 6.702897242e-16 wuc = 1.809243293e-16 puc = -3.881559468e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = -3.617169497e-01 la0 = 4.741572133e-06 wa0 = 1.195782565e-06 pa0 = -3.792236058e-12
+ ags = -5.238562694e-01 lags = 2.569241224e-06 wags = 5.157304550e-07 pags = -1.378375600e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -8.057683483e-08 lb0 = 6.589646768e-14 wb0 = 5.610419971e-14 pb0 = -4.588252431e-20
+ b1 = 7.607003178e-08 lb1 = -1.456635080e-12 wb1 = -5.296619387e-14 pb1 = 1.014228786e-18
+ keta = 2.142250194e-01 lketa = -6.253648954e-07 wketa = -1.295667662e-07 pketa = 3.845417587e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.578301750e+00 lpclm = 8.857007879e-06 wpclm = 2.846273593e-06 ppclm = -6.101515171e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -5.715063365e-03 lpdiblc2 = -3.307762063e-09 wpdiblc2 = 4.964995469e-09 ppdiblc2 = 7.643539485e-15
+ pdiblcb = 5.820108933e-02 lpdiblcb = -3.308188465e-07 wpdiblcb = -5.793142088e-08 ppdiblcb = 2.303432081e-13
+ drout = 0.56
+ pscbe1 = 1.146799543e+09 lpscbe1 = -6.853230616e+02 wpscbe1 = -3.172880548e+02 ppscbe1 = 6.270043475e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.449986400e-01 lkt1 = 1.061567109e-06 wkt1 = 1.735711697e-07 pkt1 = -7.335970491e-13
+ kt2 = -8.362615554e-02 lkt2 = 5.371792324e-07 wkt2 = 4.175183485e-08 pkt2 = -3.658229013e-13
+ at = 1.562757189e+05 lat = -6.471447193e-02 wat = 8.481160017e-03 pat = -3.372224567e-8
+ ute = -7.581647527e+00 lute = 3.155890056e-05 wute = 4.067003215e-06 pute = -2.016019040e-11
+ ua1 = -1.963254543e-08 lua1 = 9.608303450e-14 wua1 = 1.320050496e-14 pua1 = -6.100538515e-20
+ ub1 = 1.634205074e-17 lub1 = -7.613519586e-23 wub1 = -1.080888982e-23 pub1 = 4.812072319e-29
+ uc1 = -1.069321342e-10 luc1 = -1.003931456e-15 wuc1 = 6.993424884e-17 puc1 = 6.663724895e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.272467988e-03 ltvoff = 1.452366429e-08 wtvoff = 2.240838100e-09 ptvoff = -1.125585907e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.85 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.623723554e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.735077868e-07 wvth0 = -1.462399977e-08 pvth0 = -9.046474098e-14
+ k1 = 6.424935211e-01 lk1 = -6.519919438e-07 wk1 = -3.088153742e-08 pk1 = 3.731756294e-13
+ k2 = 3.093513475e-02 lk2 = 1.404631885e-07 wk2 = -5.890613301e-08 pk2 = -7.123667901e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.846493088e+00 ldsub = -4.477041017e-06 wdsub = -2.780708202e-06 pdsub = 2.714349382e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-4.404695139e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 4.744387905e-08 wvoff = 1.619807478e-07 pvoff = -6.102852672e-14
+ nfactor = 1.852926177e+00 lnfactor = -2.961415355e-06 wnfactor = 7.110895333e-07 pnfactor = 1.226866015e-12
+ eta0 = 1.213937514e+00 leta0 = -1.182496888e-06 weta0 = -7.368874447e-07 peta0 = 7.193021338e-13
+ etab = -9.811641583e-01 letab = 8.753881819e-07 wetab = 6.441974002e-07 petab = -6.288242734e-13
+ u0 = 6.755363504e-03 lu0 = 8.807252291e-09 wu0 = 1.550347924e-08 pu0 = -9.149338892e-15
+ ua = -9.031842606e-09 lua = 5.765087721e-15 wua = 5.642840652e-15 pua = -4.329117186e-21
+ ub = 1.335822209e-17 lub = -9.053194994e-24 wub = -8.061579233e-24 pub = 6.514881860e-30
+ uc = -1.187470309e-10 luc = 3.855408074e-16 wuc = 1.094374606e-16 puc = -2.468881719e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.694418099e+04 lvsat = 1.048455140e-01 wvsat = 3.014515251e-02 pvsat = -5.957092110e-8
+ a0 = 7.202927904e+00 la0 = -1.020719489e-05 wa0 = -4.065030723e-06 pa0 = 6.603846470e-12
+ ags = 4.627163445e+00 lags = -7.609874270e-06 wags = -2.974300326e-06 pags = 5.518399868e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.785220973e-07 lb0 = -1.038959060e-12 wb0 = -3.331863230e-13 pb0 = 7.234084920e-19
+ b1 = -1.260590771e-06 lb1 = 1.184788453e-12 wb1 = 8.777266633e-13 pb1 = -8.249468737e-19
+ keta = -6.862209452e-01 lketa = 1.154038791e-06 wketa = 4.591519098e-07 pketa = -7.788464108e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.310888861e+00 lpclm = -2.780833698e-06 wpclm = -1.310324341e-06 ppclm = 2.112487645e-12
+ pdiblc1 = 5.430714416e-01 lpdiblc1 = -3.024899864e-07 wpdiblc1 = -7.171716755e-08 ppdiblc1 = 1.417228766e-13
+ pdiblc2 = -2.758207008e-02 lpdiblc2 = 3.990441711e-08 wpdiblc2 = 2.254657805e-08 ppdiblc2 = -2.710005880e-14
+ pdiblcb = 1.557888629e-01 lpdiblcb = -5.236655591e-07 wpdiblcb = -1.093148461e-07 ppdiblcb = 3.318838444e-13
+ drout = 4.153991572e+00 ldrout = -7.102216130e-06 wdrout = -2.391849865e-06 pdrout = 4.726620624e-12
+ pscbe1 = 3.653269851e+08 lpscbe1 = 8.589729929e+02 wpscbe1 = 3.026549961e+02 ppscbe1 = -5.980874334e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.613969708e-05 lalpha0 = -7.135767235e-11 walpha0 = -2.514171650e-11 palpha0 = 4.968345108e-17
+ alpha1 = 2.005432075e+00 lalpha1 = -2.283290919e-06 walpha1 = -7.005176692e-07 palpha1 = 1.384318185e-12
+ beta0 = 3.755885028e+01 lbeta0 = -4.683215121e-05 wbeta0 = -1.650108287e-05 pbeta0 = 3.260838391e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.166165634e-01 lkt1 = -2.458745130e-07 wkt1 = -3.081050418e-07 pkt1 = 2.182606528e-13
+ kt2 = 4.671301857e-01 lkt2 = -5.511902008e-07 wkt2 = -3.249848058e-07 pkt2 = 3.588985769e-13
+ at = 9.019482680e+03 lat = 2.262838777e-01 wat = 8.846774109e-02 pat = -1.917866080e-7
+ ute = 1.741548466e+01 lute = -1.783883224e-05 wute = -1.199591092e-05 pute = 1.158231248e-11
+ ua1 = 5.630177954e-08 lua1 = -5.397351870e-14 wua1 = -3.508084813e-14 pua1 = 3.440513481e-20
+ ub1 = -4.245147974e-17 lub1 = 4.004881629e-23 wub1 = 2.631512563e-23 pub1 = -2.524138019e-29
+ uc1 = -1.081824386e-09 luc1 = 9.225882190e-16 wuc1 = 6.994086697e-16 puc1 = -5.775545747e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 9.036082005e-03 ltvoff = -9.799704456e-09 wtvoff = -6.700832482e-09 ptvoff = 6.414098067e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.86 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {9.087298667e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.645842488e-07 wvth0 = -2.094795072e-07 pvth0 = 9.974073466e-14
+ k1 = -5.019757873e-01 lk1 = 4.651657491e-07 wk1 = 6.860620979e-07 pk1 = -3.266588630e-13
+ k2 = 3.534422085e-01 lk2 = -1.743475764e-07 wk2 = -2.574741521e-07 pk2 = 1.225927129e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.282475902e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.307408194e-07 wvoff = 1.941734251e-07 pvoff = -9.245295793e-14
+ nfactor = -5.486117664e+00 lnfactor = 4.202489544e-06 wnfactor = 3.841972216e-06 pnfactor = -1.829301283e-12
+ eta0 = -4.616708363e-01 leta0 = 4.531247453e-07 weta0 = -4.578546857e-13 peta0 = 2.180010989e-19
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 7.428819227e-03 lu0 = 8.149867916e-09 wu0 = 1.196833064e-08 pu0 = -5.698553079e-15
+ ua = -4.719923498e-09 lua = 1.556068250e-15 wua = 2.358125433e-15 pua = -1.122788411e-21
+ ub = 6.166566058e-18 lub = -2.033160645e-24 wub = -2.708631692e-24 pub = 1.289677060e-30
+ uc = 4.892255971e-10 luc = -2.079231619e-16 wuc = -2.801246538e-16 puc = 1.333774322e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.077054884e+04 lvsat = 6.206501854e-02 wvsat = -6.029030502e-02 pvsat = 2.870638467e-8
+ a0 = -7.670831126e+00 la0 = 4.311616755e-06 wa0 = 5.271647281e-06 pa0 = -2.510021050e-12
+ ags = -6.335059408e+00 lags = 3.090746097e-06 wags = 5.230156489e-06 pags = -2.490265790e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.143712827e-06 lb0 = 5.445628508e-13 wb0 = 7.963466549e-13 pb0 = -3.791693109e-19
+ b1 = -9.143915996e-08 lb1 = 4.353747587e-14 wb1 = 6.366744118e-14 pb1 = -3.031436077e-20
+ keta = 9.751614542e-01 lketa = -4.676963786e-07 wketa = -6.613034043e-07 pketa = 3.148703577e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -1.480429790e+00 lpclm = 9.200089246e-07 wpclm = 1.666865769e-06 ppclm = -7.936547997e-13
+ pdiblc1 = 4.237879451e-01 lpdiblc1 = -1.860530712e-07 wpdiblc1 = 1.434343351e-07 ppdiblc1 = -6.829425058e-14
+ pdiblc2 = 2.591690982e-02 lpdiblc2 = -1.231786313e-08 wpdiblc2 = -1.018306457e-08 ppdiblc2 = 4.848523631e-15
+ pdiblcb = -6.530989907e-01 lpdiblcb = 2.659189948e-07 wpdiblcb = 4.503553757e-07 ppdiblcb = -2.144304072e-13
+ drout = -7.046982730e+00 ldrout = 3.831458121e-06 wdrout = 4.783699729e-06 pdrout = -2.277691654e-12
+ pscbe1 = 2.015071226e+09 lpscbe1 = -7.514017517e+02 wpscbe1 = -6.053099923e+02 ppscbe1 = 2.882098785e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -7.587468680e-05 lalpha0 = 3.798360027e-11 walpha0 = 5.028343301e-11 palpha0 = -2.394175266e-17
+ alpha1 = -1.460864150e+00 lalpha1 = 1.100285613e-06 walpha1 = 1.401035338e-06 palpha1 = -6.670833619e-13
+ beta0 = -3.749724754e+01 lbeta0 = 2.643280790e-05 wbeta0 = 3.300216575e-05 pbeta0 = -1.571351919e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = 1.554099991e-03 lkt1 = -1.335579002e-07 wkt1 = -1.649835406e-07 pkt1 = 7.855460309e-14
+ kt2 = -1.554491249e-01 lkt2 = 5.653187723e-08 wkt2 = 8.333841687e-08 pkt2 = -3.968042045e-14
+ at = 4.600295332e+05 lat = -2.139632689e-01 wat = -2.108601223e-01 pat = 1.003980952e-7
+ ute = -4.301595081e-01 lute = -4.190565268e-07 wute = -2.546560291e-07 pute = 1.212509031e-13
+ ua1 = 1.177374702e-09 lua1 = -1.646026586e-16 wua1 = 3.229120899e-16 pua1 = -1.537500708e-22
+ ub1 = -2.177482010e-18 lub1 = 7.359172347e-25 wub1 = 8.915225567e-25 pub1 = -4.244859841e-31
+ uc1 = -2.723054692e-10 luc1 = 1.323876614e-16 wuc1 = 2.103268131e-16 puc1 = -1.001441675e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.958519023e-03 ltvoff = 9.325214136e-10 wtvoff = -2.536514959e-10 ptvoff = 1.207726087e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.87 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.069956548e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.091772808e-8
+ k1 = 8.414013965e-02 lk1 = 1.860948561e-7
+ k2 = 1.045496918e-01 lk2 = -5.584088905e-08 wk2 = -1.387778781e-23 pk2 = 2.081668171e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425678e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-1.121188879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.500663643e-8
+ nfactor = 3.435621945e+00 lnfactor = -4.547186666e-8
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = 1.040834086e-23 petab = -1.301042607e-30
+ u0 = 2.128959387e-02 lu0 = 1.550254118e-9
+ ua = -1.703807103e-09 lua = 1.199866544e-16
+ ub = 1.993090002e-18 lub = -4.601845034e-26
+ uc = 1.633443546e-11 luc = 1.723734427e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.073063673e+05 lvsat = -2.944599905e-3
+ a0 = 1.280215623e+00 la0 = 4.970115974e-8
+ ags = -8.330949981e-01 lags = 4.710627705e-07 pags = -5.551115123e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.484793983e-17 lb0 = -7.880373722e-24
+ b1 = -2.675520754e-18 lb1 = 6.050315613e-25
+ keta = 6.166340678e-02 lketa = -3.274707228e-08 wketa = -1.387778781e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949620e-01 lpclm = -9.183947440e-8
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 wpdiblc1 = -5.551115123e-23 ppdiblc1 = -2.775557562e-29
+ pdiblc2 = -7.515255686e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 1.843143693e-24 ppdiblc2 = 3.117081246e-31
+ pdiblcb = -8.674421607e-02 lpdiblcb = -3.742902200e-9
+ drout = 1.449262699e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107030e+08 lpscbe1 = 1.526664888e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183450e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126009e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532619e+03 lat = 7.780439653e-3
+ ute = -1.302351205e+00 lute = -3.774660934e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591219e-16 wua1 = -8.271806126e-31
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25 wub1 = 7.703719778e-40
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = -1.292469707e-32 puc1 = 1.615587134e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.88 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820277676e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033728658e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217056813e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944838817e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083471173e-16
+ ags = 1.250000000e+00 lags = 4.460787295e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566857920e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563461134e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889157719e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866340637e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.132038907e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135939962e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034206331e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393363028e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.89 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.5e-07 wmax = 7.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-1.077060979e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 9.323666936e-08 wvth0 = 4.729775370e-07 pvth0 = -7.384882071e-14
+ k1 = 0.90707349
+ k2 = -1.811160616e-01 lk2 = 6.770416191e-09 wk2 = 5.995319769e-09 pk2 = -9.360852474e-16
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999998e-03 lcdscd = 3.262303622e-19 wcdscd = 2.012161271e-18 pcdscd = -3.141705646e-25
+ cit = 0.0
+ voff = {1.694554462e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.969838595e-07 wvoff = -1.153199572e-06 pvoff = 1.800559683e-13
+ nfactor = 2.011566944e+01 lnfactor = -2.669774261e-06 wnfactor = -1.040382246e-05 pnfactor = 1.624411224e-12
+ eta0 = 1.167676555e-09 leta0 = -1.472888359e-16 weta0 = -6.513119562e-20 peta0 = 1.016932436e-26
+ etab = -0.043998
+ u0 = 1.175812733e-01 lu0 = -1.353652246e-08 wu0 = -4.877379815e-08 pu0 = 7.615345748e-15
+ ua = -1.167043358e-09 lua = -2.205575086e-18 wua = -8.564331521e-18 pua = 1.337200466e-24
+ ub = -6.524880699e-20 lub = 3.242009357e-25 wub = 1.258884510e-24 pub = -1.965571919e-31
+ uc = 7.700399986e-11 luc = 1.717288990e-26 wuc = -1.381391623e-28 puc = 2.155839471e-35
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.864703682e+05 lvsat = -2.938539115e-02 wvsat = -8.170612732e-02 pvsat = 1.275726790e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.226508446e-18 wketa = 7.893685705e-20 pketa = -1.232347557e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.083066820e+00 lpclm = -1.411003228e-07 wpclm = -5.478978956e-07 ppclm = 8.554658583e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.058713578e-24 walpha0 = -1.577598864e-25 palpha0 = 2.463012992e-32
+ alpha1 = 0.85
+ beta0 = 1.057036139e+01 lbeta0 = 5.141203221e-07 wbeta0 = 1.996348684e-06 pbeta0 = -3.117018981e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.697880826e-02 lkt1 = -2.570601627e-08 wkt1 = -9.981743435e-08 pkt1 = 1.558509493e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.012865687e-11 wat = -3.352761269e-14 pat = 5.267793313e-21
+ ute = -2.138952857e+00 lute = 1.285300811e-07 wute = 4.990871718e-07 pute = -7.792547465e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.559757939e-02 ltvoff = -8.680783655e-09 wtvoff = -3.370781163e-08 ptvoff = 5.263002876e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.90 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.91 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-07 wk2 = -4.440892099e-22
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-07 wvoff = 1.776356839e-21
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24 wub = -1.232595164e-38
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15 pb0 = -5.293955920e-35
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13 pb1 = 1.694065895e-33
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-07 wkt2 = 2.220446049e-22
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16 puc1 = 3.308722450e-36
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.92 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-07 pk2 = 8.881784197e-28
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15 wua = -6.617444900e-30
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = -1.654361225e-30 pb0 = 3.308722450e-35
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = -8.881784197e-22 ppclm = 1.065814104e-26
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-08 ppdiblc2 = -5.551115123e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 wtvoff = -1.734723476e-24 ptvoff = -1.040834086e-29
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.93 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-6
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13 pb1 = 8.470329473e-34
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24 pub1 = -1.232595164e-44
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-09 ptvoff = -1.387778781e-29
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.94 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 peta0 = -6.938893904e-30
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = 1.318389842e-22 petab = -3.538835891e-28
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17 wuc = -4.135903063e-31
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = 1.058791184e-28 pb0 = -2.117582368e-34
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 wketa = -5.551115123e-23 pketa = 2.220446049e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = 6.776263578e-27 palpha0 = 9.317362420e-33
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-02 wat = -9.313225746e-16
+ ute = -2.370540520e+00 lute = 1.265004727e-6
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 pua1 = 3.308722450e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = -3.081487911e-39 pub1 = 3.081487911e-45
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10 wtvoff = -1.387778781e-23
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.95 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.632148963e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -7.213288526e-11
+ k1 = 6.296133048e-01 lk1 = -7.362455486e-8
+ k2 = -7.123500794e-02 lk2 = 2.785653473e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.079784331e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.824914399e-8
+ nfactor = 8.508216088e-01 lnfactor = 1.185244626e-6
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 1.193489751e-21 peta0 = 5.412337245e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.716935357e-02 lu0 = -1.249311144e-9
+ ua = -8.304373629e-10 lua = -2.958561203e-16
+ ub = 1.698955783e-18 lub = 9.402944022e-26
+ uc = 2.718870036e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.867212802e+04 lvsat = 1.094132569e-1
+ a0 = 1.024210589e+00 la0 = 1.715943729e-7
+ ags = 2.291547499e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805318e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954251e-15
+ keta = -1.155907112e-01 lketa = 5.164999443e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432982e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988834e-03 lpdiblc2 = -4.320720496e-09 ppdiblc2 = 2.775557562e-29
+ pdiblcb = 8.971602891e-02 lpdiblcb = -8.776197740e-08 wpdiblcb = 1.647987302e-22 ppdiblcb = -2.203098814e-28
+ drout = 8.432395257e-01 ldrout = 7.463925758e-8
+ pscbe1 = 1.016674453e+09 lpscbe1 = -2.760291058e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12 walpha0 = 5.421010862e-26
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690257e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136186e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908083e-9
+ at = 1.122373799e+05 lat = -4.836690423e-2
+ ute = -8.501885195e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976372e-16
+ ub1 = -7.070069559e-19 lub1 = 3.577112441e-26
+ uc1 = 7.460704527e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.376891160e-03 ltvoff = 1.131723449e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.96 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.069956548e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.091772808e-8
+ k1 = 8.414013965e-02 lk1 = 1.860948561e-7
+ k2 = 1.045496918e-01 lk2 = -5.584088905e-08 pk2 = -2.775557562e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425678e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-1.121188879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.500663643e-8
+ nfactor = 3.435621945e+00 lnfactor = -4.547186666e-8
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = -7.632783294e-23 petab = -4.510281038e-29
+ u0 = 2.128959387e-02 lu0 = 1.550254118e-9
+ ua = -1.703807103e-09 lua = 1.199866544e-16
+ ub = 1.993090002e-18 lub = -4.601845034e-26
+ uc = 1.633443546e-11 luc = 1.723734427e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.073063673e+05 lvsat = -2.944599905e-3
+ a0 = 1.280215623e+00 la0 = 4.970115974e-8
+ ags = -8.330949981e-01 lags = 4.710627705e-07 wags = 1.776356839e-21 pags = 1.332267630e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.484793983e-17 lb0 = -7.880373722e-24
+ b1 = -2.675520754e-18 lb1 = 6.050315613e-25
+ keta = 6.166340678e-02 lketa = -3.274707228e-08 wketa = 1.665334537e-22 pketa = 4.163336342e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949620e-01 lpclm = -9.183947440e-08 wpclm = 3.552713679e-21
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 wpdiblc1 = -4.440892099e-22 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -7.515255686e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 4.336808690e-25 ppdiblc2 = 8.456776945e-30
+ pdiblcb = -8.674421607e-02 lpdiblcb = -3.742902200e-9
+ drout = 1.449262699e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107030e+08 lpscbe1 = 1.526664888e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183450e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126009e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532619e+03 lat = 7.780439653e-03 pat = -2.910383046e-23
+ ute = -1.302351205e+00 lute = -3.774660934e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591219e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25 wub1 = 6.162975822e-39
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = -2.584939414e-31 puc1 = 5.169878828e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.97 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820144449e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033839681e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217143549e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944977595e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083524464e-16
+ ags = 1.250000000e+00 lags = 4.461497838e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566924534e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.562906023e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831512802e-18
+ drout = 5.033266588e-01 ldrout = 1.889137735e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866149902e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.132094418e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135939574e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034217886e-34
+ uc1 = 1.471862500e-10 luc1 = -4.392329053e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.98 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.4e-07 wmax = 6.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.807478950e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -9.864726632e-07 wvth0 = -3.719574684e-06 pvth0 = 5.807595129e-13
+ k1 = 0.90707349
+ k2 = -8.520167857e-01 lk2 = 1.115221717e-07 wk2 = 4.127503526e-07 pk2 = -6.444518905e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.45863
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000024e-03 lcdscd = -3.677003146e-18 wcdscd = -1.353256396e-17 pcdscd = 2.112914010e-24
+ cit = 0.0
+ voff = {-1.872588144e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.891381321e-06 wvoff = 1.122734315e-05 pvoff = -1.752992450e-12
+ nfactor = -1.030236525e+02 lnfactor = 1.655670690e-05 wnfactor = 6.425333190e-05 pnfactor = -1.003225823e-11
+ eta0 = 1.166700809e-09 leta0 = -1.471364686e-16 weta0 = 5.265167660e-19 peta0 = -8.220822178e-26
+ etab = -0.043998
+ u0 = -4.343177637e-01 lu0 = 7.263478558e-08 wu0 = 2.858326538e-07 pu0 = -4.462876723e-14
+ ua = -1.167043295e-09 lua = -2.205584809e-18 wua = -8.564369276e-18 pua = 1.337206361e-24
+ ub = -6.524872088e-20 lub = 3.242009223e-25 wub = 1.258884458e-24 pub = -1.965571837e-31
+ uc = 7.700399986e-11 luc = 1.744689348e-26 wuc = 9.280966473e-28 puc = -1.449634023e-34
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.502770248e+06 lvsat = 4.217290817e-01 wvsat = 1.669988452e+00 pvsat = -2.607453169e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.068967799e-18 wketa = -5.320188734e-19 pketa = 8.304468224e-26
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.083066832e+00 lpclm = -1.411003247e-07 wpclm = -5.478979030e-07 ppclm = 8.554658699e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000001e-08 lalpha0 = -1.744040838e-24 walpha0 = 1.064720415e-24 palpha0 = -1.662302159e-31
+ alpha1 = 0.85
+ beta0 = 1.057036138e+01 lbeta0 = 5.141203238e-07 wbeta0 = 1.996348691e-06 pbeta0 = -3.117018992e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -6.697881003e-02 lkt1 = -2.570601599e-08 wkt1 = -9.981743328e-08 pkt1 = 1.558509476e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.019611955e-11 wat = 2.272427082e-13 pat = -3.562308848e-20
+ ute = -2.138952848e+00 lute = 1.285300797e-07 wute = 4.990871664e-07 pute = -7.792547381e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.159933142e-01 ltvoff = 4.933793210e-08 wtvoff = 1.915810585e-07 ptvoff = -2.991270015e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.99 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.100 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.101 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = 2.067951531e-30 pb0 = -1.323488980e-35
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13 wb1 = 2.117582368e-28
+ keta = -1.746390476e-02 lketa = 8.039550078e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = 2.220446049e-22 ppclm = -5.329070518e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15 wua1 = -3.308722450e-30
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 wuc1 = 5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 wtvoff = 8.673617380e-25 ptvoff = -1.734723476e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.102 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-06 wa0 = 3.552713679e-21
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-09 ptvoff = 3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.103 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 peta0 = -1.734723476e-30
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = -3.122502257e-23 petab = -3.989863995e-29
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-06 pags = 1.776356839e-27
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = -2.646977960e-29
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = 2.646977960e-27 palpha0 = 5.505714157e-33
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-07 wkt1 = 8.881784197e-22
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-2
+ ute = -2.370540520e+00 lute = 1.265004727e-6
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = 1.240770919e-30 pua1 = 3.308722450e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = -3.851859889e-40 pub1 = 7.703719778e-46
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.104 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.632148963e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -7.213288526e-11
+ k1 = 6.296133048e-01 lk1 = -7.362455486e-8
+ k2 = -7.123500794e-02 lk2 = 2.785653473e-08 pk2 = -5.551115123e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.079784331e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.824914399e-8
+ nfactor = 8.508216088e-01 lnfactor = 1.185244626e-6
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 4.232725281e-22 peta0 = 2.081668171e-29
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.716935357e-02 lu0 = -1.249311144e-9
+ ua = -8.304373629e-10 lua = -2.958561203e-16
+ ub = 1.698955783e-18 lub = 9.402944022e-26
+ uc = 2.718870036e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.867212802e+04 lvsat = 1.094132569e-1
+ a0 = 1.024210589e+00 la0 = 1.715943729e-7
+ ags = 2.291547499e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805318e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954251e-15
+ keta = -1.155907112e-01 lketa = 5.164999443e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432982e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988834e-03 lpdiblc2 = -4.320720496e-9
+ pdiblcb = 8.971602891e-02 lpdiblcb = -8.776197740e-08 wpdiblcb = 4.770489559e-23 ppdiblcb = -1.951563910e-29
+ drout = 8.432395257e-01 ldrout = 7.463925758e-8
+ pscbe1 = 1.016674453e+09 lpscbe1 = -2.760291058e+02 wpscbe1 = -1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12 walpha0 = -1.355252716e-26
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690257e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136186e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908083e-9
+ at = 1.122373799e+05 lat = -4.836690423e-2
+ ute = -8.501885195e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976372e-16
+ ub1 = -7.070069559e-19 lub1 = 3.577112441e-26
+ uc1 = 7.460704527e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.376891160e-03 ltvoff = 1.131723449e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.105 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.069956548e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.091772808e-8
+ k1 = 8.414013965e-02 lk1 = 1.860948561e-7
+ k2 = 1.045496918e-01 lk2 = -5.584088905e-08 wk2 = 5.551115123e-23 pk2 = -3.469446952e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425678e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-1.121188879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.500663643e-8
+ nfactor = 3.435621945e+00 lnfactor = -4.547186666e-8
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = -3.469446952e-24 petab = -3.035766083e-30
+ u0 = 2.128959387e-02 lu0 = 1.550254118e-9
+ ua = -1.703807103e-09 lua = 1.199866544e-16
+ ub = 1.993090002e-18 lub = -4.601845034e-26
+ uc = 1.633443546e-11 luc = 1.723734427e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.073063673e+05 lvsat = -2.944599905e-3
+ a0 = 1.280215623e+00 la0 = 4.970115974e-8
+ ags = -8.330949981e-01 lags = 4.710627705e-07 wags = -8.881784197e-22 pags = 1.110223025e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.484793983e-17 lb0 = -7.880373722e-24
+ b1 = -2.675520754e-18 lb1 = 6.050315613e-25
+ keta = 6.166340678e-02 lketa = -3.274707228e-08 wketa = 2.775557562e-23 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949620e-01 lpclm = -9.183947440e-8
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -7.515255686e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = -4.878909776e-31
+ pdiblcb = -8.674421607e-02 lpdiblcb = -3.742902200e-9
+ drout = 1.449262699e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107030e+08 lpscbe1 = 1.526664888e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183450e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126009e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532619e+03 lat = 7.780439653e-03 pat = 7.275957614e-24
+ ute = -1.302351205e+00 lute = -3.774660934e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591219e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25 pub1 = 3.851859889e-46
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = -1.033975766e-31 puc1 = 4.523643975e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.106 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820144449e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033750863e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217074161e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944811062e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083488937e-16
+ ags = 1.250000000e+00 lags = 4.460964931e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566880125e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563599912e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889164380e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866340637e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.132038907e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135939574e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034202479e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393156233e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.107 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.1e-07 wmax = 6.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-2.146331313e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.115394559e-07 wvth0 = 1.619421207e-06 pvth0 = -2.528499495e-13
+ k1 = 0.90707349
+ k2 = 2.465068119e-02 lk2 = -2.535717996e-08 wk2 = -1.099906779e-07 pk2 = 1.717350449e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585131626e-01 ldsub = 1.824252398e-11 wdsub = 6.966803737e-11 pdsub = -1.087768868e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335147271e-19
+ cit = 0.0
+ voff = {5.965253814e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.637937736e-07 wvoff = -3.495536364e-06 pvoff = 5.457790657e-13
+ nfactor = 3.738241829e+01 lnfactor = -5.365735359e-06 wnfactor = -1.946828078e-05 pnfactor = 3.039699488e-12
+ eta0 = 1.641780072e-02 leta0 = -2.563409442e-09 weta0 = -9.789637375e-09 peta0 = 1.528514821e-15
+ etab = -0.043998
+ u0 = -8.993815695e-02 lu0 = 1.886473130e-08 wu0 = 8.048529314e-08 pu0 = -1.256665173e-14
+ ua = -1.067214444e-09 lua = -1.779246228e-17 wua = -6.809051619e-17 pua = 1.063138084e-23
+ ub = 7.948211664e-18 lub = -9.269887284e-25 wub = -3.519397727e-24 pub = 5.495046835e-31
+ uc = 3.253499464e-10 luc = -3.877574270e-17 wuc = -1.480842177e-16 puc = 2.312127742e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.779076767e+06 lvsat = -2.468213839e-01 wvsat = -8.831998500e-01 pvsat = 1.378992918e-7
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.208467322e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.993692896e-01 lpclm = 7.474772162e-08 wpclm = 2.764238727e-07 ppclm = -4.315971778e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.022661738e-24
+ alpha1 = 0.85
+ beta0 = 1.391835560e+01 lbeta0 = -8.622102004e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.708984644e-01 lkt1 = 3.736038317e-08 wkt1 = 1.410325861e-07 pkt1 = -2.202026386e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.013639849e-11
+ ute = 2.117733343e-01 lute = -2.385029035e-07 wute = -9.026085430e-07 pute = 1.409296875e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.053311047e-01 ltvoff = -1.644597737e-08 wtvoff = -5.964710865e-08 ptvoff = 9.313060956e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.108 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.109 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13 pb1 = -1.694065895e-33
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-07 wkt2 = 2.220446049e-22
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-06 wute = 7.105427358e-21
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.110 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15 wua = -6.617444900e-30
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = 3.308722450e-30 pb0 = -1.191140082e-34
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-08 wketa = -5.551115123e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = -8.881784197e-22 ppclm = 5.329070518e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 wuc1 = -2.067951531e-31 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 wtvoff = -8.673617380e-25 ptvoff = 3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.111 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-6
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.112 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 peta0 = -6.938893904e-30
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = 1.387778781e-23 petab = -2.081668171e-29
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15 pua = -3.308722450e-36
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = 1.588186776e-28 pb0 = -1.588186776e-34
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = 7.623296525e-27 palpha0 = -2.159934015e-32
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-2
+ ute = -2.370540520e+00 lute = 1.265004727e-06 wute = 1.421085472e-20
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = 1.654361225e-30 pua1 = -4.963083675e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = 1.540743956e-39 pub1 = 1.540743956e-45
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17 wuc1 = 4.135903063e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.113 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.632148963e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -7.213288526e-11
+ k1 = 6.296133048e-01 lk1 = -7.362455486e-8
+ k2 = -7.123500794e-02 lk2 = 2.785653473e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.079784331e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.824914399e-08 wvoff = -1.776356839e-21
+ nfactor = 8.508216088e-01 lnfactor = 1.185244626e-6
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 3.885780586e-22 peta0 = -3.885780586e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.716935357e-02 lu0 = -1.249311144e-9
+ ua = -8.304373629e-10 lua = -2.958561203e-16
+ ub = 1.698955783e-18 lub = 9.402944022e-26
+ uc = 2.718870036e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -2.867212802e+04 lvsat = 1.094132569e-1
+ a0 = 1.024210589e+00 la0 = 1.715943729e-7
+ ags = 2.291547499e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805318e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954251e-15
+ keta = -1.155907112e-01 lketa = 5.164999443e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432982e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988834e-03 lpdiblc2 = -4.320720496e-9
+ pdiblcb = 8.971602891e-02 lpdiblcb = -8.776197740e-08 wpdiblcb = 6.765421556e-23 ppdiblcb = 7.632783294e-29
+ drout = 8.432395257e-01 ldrout = 7.463925758e-8
+ pscbe1 = 1.016674453e+09 lpscbe1 = -2.760291058e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690257e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136186e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908083e-9
+ at = 1.122373799e+05 lat = -4.836690423e-2
+ ute = -8.501885195e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976372e-16
+ ub1 = -7.070069559e-19 lub1 = 3.577112441e-26
+ uc1 = 7.460704527e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.376891160e-03 ltvoff = 1.131723449e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.114 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.069956548e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.091772808e-8
+ k1 = 8.414013965e-02 lk1 = 1.860948561e-7
+ k2 = 1.045496918e-01 lk2 = -5.584088905e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425678e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-1.121188879e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.500663643e-8
+ nfactor = 3.435621945e+00 lnfactor = -4.547186666e-8
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = 6.245004514e-23 petab = 5.204170428e-30
+ u0 = 2.128959387e-02 lu0 = 1.550254118e-9
+ ua = -1.703807103e-09 lua = 1.199866544e-16
+ ub = 1.993090002e-18 lub = -4.601845034e-26
+ uc = 1.633443546e-11 luc = 1.723734427e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.073063673e+05 lvsat = -2.944599905e-3
+ a0 = 1.280215623e+00 la0 = 4.970115974e-8
+ ags = -8.330949981e-01 lags = 4.710627705e-07 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 3.484793983e-17 lb0 = -7.880373722e-24
+ b1 = -2.675520754e-18 lb1 = 6.050315613e-25
+ keta = 6.166340678e-02 lketa = -3.274707228e-08 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949620e-01 lpclm = -9.183947440e-8
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 ppdiblc1 = 1.110223025e-28
+ pdiblc2 = -7.515255686e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 1.214306433e-23 ppdiblc2 = -3.252606517e-31
+ pdiblcb = -8.674421607e-02 lpdiblcb = -3.742902200e-9
+ drout = 1.449262699e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107030e+08 lpscbe1 = 1.526664888e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183450e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126009e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532619e+03 lat = 7.780439653e-3
+ ute = -1.302351205e+00 lute = -3.774660934e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591219e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = 1.550963649e-31 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.115 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820499721e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033662045e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217074161e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944977595e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083453410e-16
+ ags = 1.250000000e+00 lags = 4.460787295e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.567102169e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563461134e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831512802e-18
+ drout = 5.033266588e-01 ldrout = 1.889155499e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866531372e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.131983396e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135940608e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034217886e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393156233e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.116 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 6.0e-07 wmax = 6.1e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {2.044786439e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.449339251e-08 wvth0 = 2.881998430e-07 pvth0 = -4.499837069e-14
+ k1 = 0.90707349
+ k2 = -7.265154737e-02 lk2 = -1.016479920e-08 wk2 = -5.489017732e-08 pk2 = 8.570332727e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585131590e-01 ldsub = 1.824309235e-11 wdsub = 6.967009877e-11 pdsub = -1.087801054e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335043187e-19
+ cit = 0.0
+ voff = {-2.075300001e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.749089762e-17
+ nfactor = 1.473935798e+01 lnfactor = -1.830338495e-06 wnfactor = -6.645923302e-06 pnfactor = 1.037667881e-12
+ eta0 = 1.641776644e-02 leta0 = -2.563404346e-09 weta0 = -9.789618892e-09 peta0 = 1.528511935e-15
+ etab = -0.043998
+ u0 = -2.357740547e-01 lu0 = 4.163496504e-08 wu0 = 1.630695370e-07 pu0 = -2.546102523e-14
+ ua = -1.067214413e-09 lua = -1.779246712e-17 wua = -6.809053374e-17 pua = 1.063138358e-23
+ ub = 7.948211668e-18 lub = -9.269887290e-25 wub = -3.519397730e-24 pub = 5.495046839e-31
+ uc = 3.253499468e-10 luc = -3.877574275e-17 wuc = -1.480842179e-16 puc = 2.312127745e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -7.905150410e+04 lvsat = 4.329933190e-02 wvsat = 1.690247437e-01 pvsat = -2.639084739e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.208189766e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.993692910e-01 lpclm = 7.474772183e-08 wpclm = 2.764238734e-07 ppclm = -4.315971790e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.022714678e-24
+ alpha1 = 0.85
+ beta0 = 1.391835560e+01 lbeta0 = -8.622102004e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.708984687e-01 lkt1 = 3.736038383e-08 wkt1 = 1.410325885e-07 pkt1 = -2.202026424e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.013628207e-11
+ ute = 2.117733753e-01 lute = -2.385029099e-07 wute = -9.026085663e-07 pute = 1.409296911e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.117 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.118 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-07 wk1 = -1.776356839e-21
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13 pb1 = -8.470329473e-34
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+03 ppscbe1 = -7.629394531e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16 wuc1 = 1.033975766e-31 puc1 = 8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.119 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 pb0 = 9.926167351e-36
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-08 wketa = -2.775557562e-23
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 wuc1 = -1.033975766e-31
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 wtvoff = -4.336808690e-25 ptvoff = 5.204170428e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.120 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-6
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-08 wpdiblcb = -1.110223025e-22
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.121 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 weta0 = 1.734723476e-24
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = -7.112366252e-23 petab = -1.457167720e-28
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = 5.293955920e-29 pb0 = 2.117582368e-34
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 pketa = -8.326672685e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = -5.082197684e-27 palpha0 = -4.658681210e-33
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-2
+ ute = -2.370540520e+00 lute = 1.265004727e-06 wute = 7.105427358e-21
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = 8.271806126e-31 pua1 = -1.654361225e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 pub1 = 7.703719778e-46
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.122 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {9.463205491e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -3.740353524e-07 wvth0 = -2.131147787e-07 pvth0 = 2.080290077e-13
+ k1 = 6.296133055e-01 lk1 = -7.362455560e-08 wk1 = -4.224496308e-16 pk1 = 4.123679176e-22
+ k2 = -7.007651624e-02 lk2 = 2.672568927e-08 wk2 = -6.444480799e-10 pk2 = 6.290689709e-16
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939289e-01 ldsub = 4.676284059e-08 wdsub = -1.245989978e-16 pdsub = 1.216262646e-22
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.427250110e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.146946522e-06 wvoff = 1.178912687e-06 pvoff = -1.150779115e-12
+ nfactor = -3.351275102e+01 lnfactor = 3.472876496e-05 wnfactor = 1.911583691e-05 pnfactor = -1.865965658e-11
+ eta0 = -4.616715920e-01 leta0 = 4.531251054e-07 weta0 = 2.850791964e-16 peta0 = -2.782767558e-22
+ etab = -1.641277801e-01 letab = 7.784955976e-08 wetab = 5.727862629e-17 petab = -5.591149765e-23
+ u0 = -4.618052436e-02 lu0 = 7.035014530e-08 wu0 = 4.080321679e-08 pu0 = -3.982948883e-14
+ ua = -8.304373597e-10 lua = -2.958561234e-16 wua = -1.795418681e-24 pua = 1.752574034e-30
+ ub = 1.698955786e-18 lub = 9.402943746e-26 wub = -1.572551074e-33 pub = 1.535024714e-39
+ uc = 2.718870047e-11 luc = 1.206923788e-17 wuc = -6.421196300e-26 puc = 6.267950752e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.355513382e+05 lvsat = 7.018099016e-01 wvsat = 3.375959808e-01 pvsat = -3.295395903e-7
+ a0 = 1.024210583e+00 la0 = 1.715943783e-07 wa0 = 3.105625979e-15 pa0 = -3.031509266e-21
+ ags = 2.291547474e+00 lags = -1.016691985e-06 wags = 1.372291081e-14 pags = -1.339542877e-20
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793340e-07 lb0 = -8.083805273e-14 wb0 = 2.598993544e-22 pb0 = -2.536971674e-28
+ b1 = 1.357375680e-08 lb1 = -6.462954286e-15 wb1 = -1.995429629e-23 pb1 = 1.947811819e-29
+ keta = -1.155907120e-01 lketa = 5.164999526e-08 wketa = 4.734999060e-16 pketa = -4.622001670e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894407e+00 lpclm = -3.890433046e-07 wpclm = -3.627615541e-15 ppclm = 3.541048343e-21
+ pdiblc1 = 6.603681741e-01 lpdiblc1 = -2.986974345e-07 wpdiblc1 = 6.799645291e-16 ppdiblc1 = -6.637375094e-22
+ pdiblc2 = 9.120988864e-03 lpdiblc2 = -4.320720524e-09 wpdiblc2 = -1.638658653e-17 ppdiblc2 = 1.599552435e-23
+ pdiblcb = 8.971602867e-02 lpdiblcb = -8.776197717e-08 wpdiblcb = 1.316537825e-16 ppdiblcb = -1.285117945e-22
+ drout = 8.432395265e-01 ldrout = 7.463925678e-08 wdrout = -4.569820078e-16 pdrout = 4.460751768e-22
+ pscbe1 = 1.016674444e+09 lpscbe1 = -2.760290966e+02 wpscbe1 = 5.261962891e-06 ppscbe1 = -5.136388779e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680628e-06 lalpha0 = -1.505866098e-12 walpha0 = 6.176455831e-21 palpha0 = -6.029058546e-27
+ alpha1 = 0.85
+ beta0 = 1.693644136e+01 lbeta0 = 5.149689774e-07 wbeta0 = -2.750090289e-14 pbeta0 = 2.684464562e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693354e-01 lkt1 = -3.990136108e-09 wkt1 = 4.413180932e-17 pkt1 = -4.307931789e-23
+ kt2 = -1.799095059e-02 lkt2 = -8.916908071e-09 wkt2 = 7.193023954e-18 pkt2 = -7.021383475e-24
+ at = 1.122373789e+05 lat = -4.836690327e-02 wat = 5.465282593e-10 pat = -5.334857851e-16
+ ute = -8.501885175e-01 lute = -2.190655954e-07 wute = -1.129670579e-15 pute = 1.102709035e-21
+ ua1 = 1.709985083e-09 lua1 = -4.181976331e-16 wua1 = 2.340299094e-24 pua1 = -2.284447859e-30
+ ub1 = -7.070069568e-19 lub1 = 3.577112531e-26 wub1 = 5.134590861e-34 pub1 = -5.012040087e-40
+ uc1 = 7.460704537e-11 luc1 = -3.278987573e-17 wuc1 = -5.686804673e-26 puc1 = 5.551085014e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.906562752e-02 ltvoff = 5.646763981e-08 wtvoff = 3.153492364e-08 ptvoff = -3.078237422e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.123 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-1.592156508e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.523502317e-07 wvth0 = 4.262295575e-07 pvth0 = -9.638584721e-14
+ k1 = 8.414013813e-02 lk1 = 1.860948564e-07 wk1 = 8.448974853e-16 pk1 = -1.910622771e-22
+ k2 = 1.022327084e-01 lk2 = -5.531693569e-08 wk2 = 1.288896160e-09 pk2 = -2.914658220e-16
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425674e-01 ldsub = 6.388057806e-08 wdsub = 2.491997719e-16 pdsub = -5.635314437e-23
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {4.126424466e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.734938763e-07 wvoff = -2.357825374e-06 pvoff = 5.331891987e-13
+ nfactor = 7.216276721e+01 lnfactor = -1.558715359e-05 wnfactor = -3.823167382e-05 pnfactor = 8.645557791e-12
+ eta0 = 9.325986808e-01 leta0 = -2.107371652e-07 weta0 = -5.701608075e-16 peta0 = 1.289333085e-22
+ etab = 3.860778713e-02 letab = -1.868014228e-08 wetab = -1.145570479e-16 petab = 2.590545660e-23
+ u0 = 1.679893497e-01 lu0 = -3.162384187e-08 wu0 = -8.160643359e-08 pu0 = 1.845415247e-14
+ ua = -1.703807110e-09 lua = 1.199866558e-16 wua = 3.590843979e-24 pua = -8.120200463e-31
+ ub = 1.993089997e-18 lub = -4.601844906e-26 wub = 3.145102147e-33 pub = -7.112212766e-40
+ uc = 1.633443523e-11 luc = 1.723734432e-17 wuc = 1.284239260e-25 puc = -2.904122563e-32
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.421064788e+06 lvsat = -2.774190740e-01 wvsat = -6.751919615e-01 pvsat = 1.526852094e-7
+ a0 = 1.280215634e+00 la0 = 4.970115722e-08 wa0 = -6.211244852e-15 pa0 = 1.404586669e-21
+ ags = -8.330949487e-01 lags = 4.710627593e-07 wags = -2.744582339e-14 pags = 6.206488878e-21
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 9.692640833e-16 lb0 = -2.191855027e-22 wb0 = -5.197988811e-22 pb0 = 1.175452398e-28
+ b1 = -7.441720181e-17 lb1 = 1.682840835e-23 wb1 = 3.990860582e-23 pb1 = -9.024772486e-30
+ keta = 6.166340848e-02 lketa = -3.274707267e-08 wketa = -9.469993401e-16 pketa = 2.141506625e-22
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949490e-01 lpclm = -9.183947145e-08 wpclm = 7.255232859e-15 ppclm = -1.640669378e-21
+ pdiblc1 = -2.599865108e-01 lpdiblc1 = 1.395165637e-07 wpdiblc1 = -1.359929169e-15 ppdiblc1 = 3.075291410e-22
+ pdiblc2 = -7.515255745e-03 lpdiblc2 = 3.600394438e-09 wpdiblc2 = 3.277315311e-17 ppdiblc2 = -7.411186628e-24
+ pdiblcb = -8.674421560e-02 lpdiblcb = -3.742902307e-09 wpdiblcb = -2.633075979e-16 ppdiblcb = 5.954337023e-23
+ drout = 1.449262698e+00 ldrout = -2.139101919e-07 wdrout = 9.139604629e-16 pdrout = -2.066791183e-22
+ pscbe1 = 1.163107219e+08 lpscbe1 = 1.526664846e+02 wpscbe1 = -1.052392387e-05 ppscbe1 = 2.379837990e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183472e-06 lalpha0 = -1.670372440e-12 walpha0 = -1.235289811e-20 palpha0 = 2.793436733e-27
+ alpha1 = 0.85
+ beta0 = 2.136300361e+01 lbeta0 = -1.592676664e-06 wbeta0 = 5.500186262e-14 pbeta0 = -1.243789427e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121571e-01 lkt1 = 1.636126006e-08 wkt1 = -8.826450681e-17 pkt1 = 1.995958954e-23
+ kt2 = -4.380991829e-02 lkt2 = 3.376431932e-09 wkt2 = -1.438626995e-17 pkt2 = 3.253203262e-24
+ at = -5.685530654e+03 lat = 7.780439208e-03 wat = -1.093056344e-09 pat = 2.471793850e-16
+ ute = -1.302351209e+00 lute = -3.774660016e-09 wute = 2.259334053e-15 pute = -5.109175305e-22
+ ua1 = 1.605522263e-09 lua1 = -3.684591238e-16 wua1 = -4.680594879e-24 pua1 = 1.058450386e-30
+ ub1 = -1.843635239e-18 lub1 = 5.769607691e-25 wub1 = -1.026915091e-33 pub1 = 2.322232401e-40
+ uc1 = -1.222035416e-10 luc1 = 6.091872993e-17 wuc1 = 1.137358867e-25 puc1 = -2.571980467e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.133774727e-01 ltvoff = -2.563872817e-08 wtvoff = -6.306984728e-08 ptvoff = 1.426236298e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.124 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820322085e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033750863e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217039466e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944755551e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083453410e-16
+ ags = 1.250000000e+00 lags = 4.460787295e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566835716e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563461134e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889155499e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866531372e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.132038907e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135940608e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034217886e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393569824e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.125 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.8e-07 wmax = 6.0e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.909930288e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.418174814e-10 wvth0 = 1.288170480e-07 pvth0 = -2.011297860e-14
+ k1 = 0.90707349
+ k2 = -6.834566699e-01 lk2 = 8.520386941e-08 wk2 = 2.848897178e-07 pk2 = -4.448154099e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585131590e-01 ldsub = 1.824309234e-11 wdsub = 6.967009872e-11 pdsub = -1.087801053e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335112576e-19
+ cit = 0.0
+ voff = {-2.075300001e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.749089762e-17
+ nfactor = -1.069954111e+01 lnfactor = 2.141589454e-06 wnfactor = 7.505278364e-06 pnfactor = -1.171844143e-12
+ eta0 = 1.641776644e-02 leta0 = -2.563404346e-09 weta0 = -9.789618892e-09 peta0 = 1.528511935e-15
+ etab = -0.043998
+ u0 = 5.288906197e-01 lu0 = -7.775671857e-08 wu0 = -2.622996574e-07 pu0 = 4.095441931e-14
+ ua = -1.067214413e-09 lua = -1.779246712e-17 wua = -6.809053374e-17 pua = 1.063138358e-23
+ ub = 7.948211668e-18 lub = -9.269887290e-25 wub = -3.519397730e-24 pub = 5.495046839e-31
+ uc = 3.253499468e-10 luc = -3.877574275e-17 wuc = -1.480842179e-16 puc = 2.312127745e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 2.394472124e+04 lvsat = 2.721791326e-02 wvsat = 1.117297975e-01 pvsat = -1.744504367e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.208467322e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.993692910e-01 lpclm = 7.474772183e-08 wpclm = 2.764238734e-07 ppclm = -4.315971790e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.022608799e-24
+ alpha1 = 0.85
+ beta0 = 1.391835560e+01 lbeta0 = -8.622102004e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.708984687e-01 lkt1 = 3.736038383e-08 wkt1 = 1.410325885e-07 pkt1 = -2.202026424e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.013628207e-11
+ ute = 2.117733753e-01 lute = -2.385029099e-07 wute = -9.026085663e-07 pute = 1.409296911e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.126 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.127 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-07 wvth0 = -8.881784197e-22
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-07 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.128 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = -3.722312756e-30 pb0 = 2.481541838e-35
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = 4.440892099e-22 ppclm = -8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 puc1 = -4.135903063e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 wtvoff = 2.168404345e-25
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.129 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-6
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-09 ptvoff = 3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.130 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-08 wk2 = 1.110223025e-22
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-9
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = 4.683753385e-23 petab = 8.326672685e-29
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15 pua = -8.271806126e-37
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 pb0 = 7.940933881e-35
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 pketa = 8.326672685e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = 7.411538288e-28 palpha0 = 6.140988868e-33
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-02 wat = 2.328306437e-16
+ ute = -2.370540520e+00 lute = 1.265004727e-6
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = 4.135903063e-31 pua1 = 8.271806126e-37
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = -7.703719778e-40 pub1 = -1.155557967e-45
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.131 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.489274262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.387438106e-8
+ k1 = 6.296133047e-01 lk1 = -7.362455483e-8
+ k2 = -7.127821251e-02 lk2 = 2.789870827e-08 wk2 = -1.110223025e-22
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.289427140e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.099533237e-9
+ nfactor = 2.132370221e+00 lnfactor = -6.572110951e-8
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = -4.163336342e-23 peta0 = -3.295974604e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.990485012e-02 lu0 = -3.919527800e-9
+ ua = -8.304373631e-10 lua = -2.958561202e-16
+ ub = 1.698955783e-18 lub = 9.402944032e-26
+ uc = 2.718870035e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.039288954e+03 lvsat = 8.732052794e-2
+ a0 = 1.024210589e+00 la0 = 1.715943727e-7
+ ags = 2.291547500e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805320e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954249e-15
+ keta = -1.155907111e-01 lketa = 5.164999439e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432980e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988833e-03 lpdiblc2 = -4.320720495e-9
+ pdiblcb = 8.971602892e-02 lpdiblcb = -8.776197741e-08 wpdiblcb = -5.377642776e-23 ppdiblcb = 4.553649124e-30
+ drout = 8.432395256e-01 ldrout = 7.463925761e-8
+ pscbe1 = 1.016674454e+09 lpscbe1 = -2.760291061e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136189e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908084e-9
+ at = 1.122373800e+05 lat = -4.836690427e-2
+ ute = -8.501885196e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976374e-16
+ ub1 = -7.070069558e-19 lub1 = 3.577112438e-26
+ uc1 = 7.460704526e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.627520928e-04 ltvoff = -9.319638031e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.132 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.355705950e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.737955077e-8
+ k1 = 8.414013971e-02 lk1 = 1.860948561e-7
+ k2 = 1.046361009e-01 lk2 = -5.586042927e-08 pk2 = 1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425679e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-2.701903262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.073900634e-8
+ nfactor = 8.725247214e-01 lnfactor = 5.341366871e-7
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = -6.938893904e-24 petab = -7.372574773e-30
+ u0 = 1.581860078e-02 lu0 = 2.787442612e-9
+ ua = -1.703807103e-09 lua = 1.199866543e-16
+ ub = 1.993090003e-18 lub = -4.601845039e-26
+ uc = 1.633443547e-11 luc = 1.723734426e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.620406891e+05 lvsat = 7.291599488e-3
+ a0 = 1.280215623e+00 la0 = 4.970115984e-8
+ ags = -8.330949999e-01 lags = 4.710627709e-07 wags = 4.440892099e-22 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.166340672e-02 lketa = -3.274707227e-08 wketa = 1.387778781e-23 pketa = 2.775557562e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949625e-01 lpclm = -9.183947451e-8
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 ppdiblc1 = -1.110223025e-28
+ pdiblc2 = -7.515255684e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 4.119968255e-24 ppdiblc2 = -2.927345866e-30
+ pdiblcb = -8.674421609e-02 lpdiblcb = -3.742902196e-9
+ drout = 1.449262700e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107023e+08 lpscbe1 = 1.526664890e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183449e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126010e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532692e+03 lat = 7.780439669e-03 pat = 7.275957614e-24
+ ute = -1.302351205e+00 lute = -3.774660968e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591218e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25 wub1 = 1.540743956e-39
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = 1.292469707e-32 puc1 = 4.846761402e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.228278134e-03 ltvoff = 9.561659042e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.133 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820144449e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033750863e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217039466e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944811062e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083453410e-16
+ ags = 1.250000000e+00 lags = 4.460964931e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566880125e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563599912e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889155499e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866245270e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.132038907e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135939832e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034202479e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393569824e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.134 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.5e-07 wmax = 5.8e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {2.010309021e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.374617392e-07 wvth0 = -6.859647707e-07 pvth0 = 1.071037954e-13
+ k1 = 0.90707349
+ k2 = -2.400899080e-01 lk2 = 1.597835667e-08 wk2 = 4.712010405e-08 pk2 = -7.357144565e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.585131559e-01 ldsub = 1.824357490e-11 wdsub = 6.967175620e-11 pdsub = -1.087826933e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335147271e-19
+ cit = 0.0
+ voff = {-5.216171058e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.820291802e-07 wvoff = 2.686044044e-06 pvoff = -4.193881728e-13
+ nfactor = -1.709154446e+01 lnfactor = 3.139611289e-06 wnfactor = 1.093319470e-05 pnfactor = -1.707065288e-12
+ eta0 = 1.641773873e-02 leta0 = -2.563400019e-09 weta0 = -9.789604030e-09 peta0 = 1.528509615e-15
+ etab = -0.043998
+ u0 = -1.745137978e-01 lu0 = 3.207003357e-08 wu0 = 1.149234704e-07 pu0 = -1.794369098e-14
+ ua = -1.067214387e-09 lua = -1.779247122e-17 wua = -6.809054781e-17 pua = 1.063138577e-23
+ ub = 7.948211672e-18 lub = -9.269887297e-25 wub = -3.519397732e-24 pub = 5.495046843e-31
+ uc = 3.253499472e-10 luc = -3.877574281e-17 wuc = -1.480842181e-16 puc = 2.312127748e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -3.917240636e+04 lvsat = 3.707276909e-02 wvsat = 1.455783769e-01 pvsat = -2.273002546e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.700000007e-02 lketa = 9.208522833e-18
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.993692922e-01 lpclm = 7.474772202e-08 wpclm = 2.764238741e-07 ppclm = -4.315971801e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000002e-08 lalpha0 = -2.022661738e-24
+ alpha1 = 0.85
+ beta0 = 1.391835560e+01 lbeta0 = -8.622102004e-9
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.708984723e-01 lkt1 = 3.736038441e-08 wkt1 = 1.410325905e-07 pkt1 = -2.202026454e-14
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.013628207e-11
+ ute = 2.117734108e-01 lute = -2.385029154e-07 wute = -9.026085853e-07 pute = 1.409296941e-13
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -9.041211588e-02 ltvoff = 1.411658612e-08 wtvoff = 4.848639033e-08 ptvoff = -7.570471040e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.135 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.136 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-07 wa0 = -7.105427358e-21
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-07 ppclm = 8.881784197e-28
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+03 ppscbe1 = -1.525878906e-17
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.137 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = -1.654361225e-30 pb0 = -3.970466940e-35
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = 4.440892099e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 wuc1 = 2.067951531e-31 puc1 = -8.271806126e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.138 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-06 wdsub = -3.552713679e-21
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-06 wa0 = -7.105427358e-21
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15 pua1 = -1.323488980e-35
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-09 ptvoff = -6.938893904e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.139 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-7
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 peta0 = -6.938893904e-30
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = -1.804112415e-22 petab = 1.179611964e-28
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15 pua = 3.308722450e-36
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = 5.293955920e-29 pb0 = 3.176373552e-34
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 wketa = 5.551115123e-23 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 palpha0 = -1.990527426e-32
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-2
+ ute = -2.370540520e+00 lute = 1.265004727e-6
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = -1.654361225e-30 pua1 = 6.617444900e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = -1.540743956e-39
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.140 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.489274262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.387438106e-8
+ k1 = 6.296133047e-01 lk1 = -7.362455483e-8
+ k2 = -7.127821251e-02 lk2 = 2.789870827e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.289427140e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.099533237e-9
+ nfactor = 2.132370221e+00 lnfactor = -6.572110951e-8
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 7.355227538e-22 peta0 = 3.469446952e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.990485012e-02 lu0 = -3.919527800e-9
+ ua = -8.304373631e-10 lua = -2.958561202e-16
+ ub = 1.698955783e-18 lub = 9.402944032e-26
+ uc = 2.718870035e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.039288954e+03 lvsat = 8.732052794e-02 pvsat = -2.328306437e-22
+ a0 = 1.024210589e+00 la0 = 1.715943727e-7
+ ags = 2.291547500e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805320e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954249e-15
+ keta = -1.155907111e-01 lketa = 5.164999439e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432980e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988833e-03 lpdiblc2 = -4.320720495e-9
+ pdiblcb = 8.971602892e-02 lpdiblcb = -8.776197741e-08 wpdiblcb = -1.249000903e-22 ppdiblcb = 4.770489559e-29
+ drout = 8.432395256e-01 ldrout = 7.463925761e-8
+ pscbe1 = 1.016674454e+09 lpscbe1 = -2.760291061e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136189e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908084e-9
+ at = 1.122373800e+05 lat = -4.836690427e-2
+ ute = -8.501885196e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976374e-16
+ ub1 = -7.070069558e-19 lub1 = 3.577112438e-26
+ uc1 = 7.460704526e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.627520928e-04 ltvoff = -9.319638031e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.141 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.355705950e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.737955077e-8
+ k1 = 8.414013971e-02 lk1 = 1.860948561e-7
+ k2 = 1.046361009e-01 lk2 = -5.586042927e-08 wk2 = -1.110223025e-22 pk2 = -8.326672685e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425679e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-09 pcdscd = -6.938893904e-30
+ cit = 0.0
+ voff = {-2.701903262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.073900634e-8
+ nfactor = 8.725247214e-01 lnfactor = 5.341366871e-7
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = -4.510281038e-23 petab = 2.428612866e-29
+ u0 = 1.581860078e-02 lu0 = 2.787442612e-9
+ ua = -1.703807103e-09 lua = 1.199866543e-16
+ ub = 1.993090003e-18 lub = -4.601845039e-26
+ uc = 1.633443547e-11 luc = 1.723734426e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.620406891e+05 lvsat = 7.291599488e-3
+ a0 = 1.280215623e+00 la0 = 4.970115984e-8
+ ags = -8.330949999e-01 lags = 4.710627709e-07 wags = 1.776356839e-21 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.166340672e-02 lketa = -3.274707227e-08 pketa = -4.163336342e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949625e-01 lpclm = -9.183947451e-08 wpclm = -3.552713679e-21
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 ppdiblc1 = -2.220446049e-28
+ pdiblc2 = -7.515255684e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = -5.204170428e-24 ppdiblc2 = 2.710505431e-30
+ pdiblcb = -8.674421609e-02 lpdiblcb = -3.742902196e-9
+ drout = 1.449262700e+00 ldrout = -2.139101923e-07 wdrout = -7.105427358e-21
+ pscbe1 = 1.163107023e+08 lpscbe1 = 1.526664890e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183449e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126010e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532692e+03 lat = 7.780439669e-03 pat = 1.455191523e-23
+ ute = -1.302351205e+00 lute = -3.774660968e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591218e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25 pub1 = 7.703719778e-46
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = 1.550963649e-31 puc1 = -3.877409121e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.228278134e-03 ltvoff = 9.561659042e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.142 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820499721e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033839681e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217004772e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944755551e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083453410e-16
+ ags = 1.250000000e+00 lags = 4.461142566e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566746898e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563738690e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831956891e-18
+ drout = 5.033266588e-01 ldrout = 1.889173262e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866531372e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.131983396e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135939574e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034217886e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393156233e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.143 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.4e-07 wmax = 5.5e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-4.661540403e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 8.042541424e-07 wvth0 = 2.691872499e-06 pvth0 = -4.202982045e-13
+ k1 = 0.90707349
+ k2 = 8.390312248e-02 lk2 = -3.460861914e-08 wk2 = -1.169117354e-07 pk2 = 1.825413072e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.467965476e+00 ldsub = -3.137296038e-07 wdsub = -1.017279868e-06 pdsub = 1.588340094e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335181965e-19
+ cit = 0.0
+ voff = {1.481839317e+01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -2.346087540e-06 wvoff = -7.457095204e-06 pvoff = 1.164321017e-12
+ nfactor = 6.899071993e+01 lnfactor = -1.030092914e-05 wnfactor = -3.264870628e-05 pnfactor = 5.097638404e-12
+ eta0 = -1.136608897e-02 leta0 = 1.774655702e-09 weta0 = 4.276847823e-09 peta0 = -6.677699117e-16
+ etab = -0.043998
+ u0 = 1.419713830e+00 lu0 = -2.168462913e-07 wu0 = -6.922052814e-07 pu0 = 1.080781638e-13
+ ua = -1.477932634e-09 lua = 4.633543300e-17 wua = 1.398487077e-16 pua = -2.183541783e-23
+ ub = 6.883165008e-18 lub = -7.606966037e-25 wub = -2.980183777e-24 pub = 4.653139742e-31
+ uc = -2.014268080e-10 luc = 4.347307263e-17 wuc = 1.186133710e-16 puc = -1.851981730e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.115674128e+06 lvsat = -1.432403494e-01 wvsat = -4.390996363e-01 pvsat = 6.855926082e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.229130883e-01 lketa = 1.242706859e-07 wketa = 4.029564701e-07 pketa = -6.291601142e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.088112420e-03 lpclm = 2.674255270e-08 wpclm = 1.207637244e-07 ppclm = -1.885556487e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.999997574e-08 lalpha0 = 3.788690917e-21 walpha0 = 1.229165593e-20 palpha0 = -1.919170088e-27
+ alpha1 = 0.85
+ beta0 = 1.391835537e+01 lbeta0 = -8.622065789e-09 wbeta0 = 1.174323643e-13 pbeta0 = -1.833538477e-20
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.923331776e-01 lkt1 = -6.133686455e-09 wkt1 = -4.101782025e-15 pkt1 = 6.404361486e-22
+ kt2 = -0.028878939
+ at = 5.372048954e+04 lat = -3.982814960e-10 wat = -1.324324869e-09 pat = 2.067746827e-16
+ ute = -1.132927112e+00 lute = -2.854675466e-08 wute = -2.218109154e-07 pute = 3.463266909e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 2.712363476e-01 ltvoff = -4.234975837e-08 wtvoff = -1.346097171e-07 ptvoff = 2.101742279e-14
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.144 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.145 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.921290502e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.208157421e-7
+ k1 = 6.123320250e-01 lk1 = -8.854283449e-7
+ k2 = -5.774281186e-02 lk2 = 3.240715930e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.541606888e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.500776891e-7
+ nfactor = 2.598709674e+00 lnfactor = 2.648900776e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.284798892e-02 lu0 = 3.954098501e-8
+ ua = -1.241809818e-09 lua = 3.755336140e-15
+ ub = 1.685065637e-18 lub = -1.765203975e-24
+ uc = 6.330548048e-11 luc = -2.950171746e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.390915283e+00 la0 = -5.656299401e-7
+ ags = 3.208651839e-01 lags = 4.797232332e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.011435769e-09 lb0 = -6.860719398e-15
+ b1 = -3.240077754e-09 lb1 = 6.604725378e-13 pb1 = -8.470329473e-34
+ keta = -2.660376772e-03 lketa = -3.767945174e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -9.712120000e-03 lpclm = 5.311079250e-7
+ pdiblc1 = 0.39
+ pdiblc2 = 5.516568119e-04 lpdiblc2 = 8.163660446e-9
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -7.410457490e+07 lpscbe1 = 5.974953667e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.832161327e-01 lkt1 = -6.320184307e-8
+ kt2 = -3.546454717e-02 lkt2 = 1.187904134e-7
+ at = 1.982637300e+05 lat = -4.647194343e-1
+ ute = -1.015897703e+00 lute = -1.987671409e-6
+ ua1 = 1.029872646e-09 lua1 = 1.820372413e-15
+ ub1 = -3.826688949e-19 lub1 = -3.731564281e-24
+ uc1 = 6.931016453e-11 luc1 = -7.089890741e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.407269502e-04 ltvoff = -3.581260738e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.146 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.232032033e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.296407051e-8
+ k1 = 4.369481614e-01 lk1 = 5.134572035e-7
+ k2 = 1.222721969e-02 lk2 = -2.340188946e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.512913721e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.271916286e-7
+ nfactor = 2.801850510e+00 lnfactor = -1.355388858e-06 wnfactor = -7.105427358e-21
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.600560204e-02 lu0 = 1.435543330e-8
+ ua = -9.768594712e-10 lua = 1.642056141e-15
+ ub = 1.627914685e-18 lub = -1.309360213e-24
+ uc = 9.599342154e-12 luc = 1.333502887e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.409463060e+00 la0 = -7.135695335e-7
+ ags = 3.609702746e-01 lags = 1.598395755e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.142758974e-09 lb0 = 7.413051884e-14 wb0 = 6.203854594e-30 pb0 = -1.158052858e-35
+ b1 = 1.158243842e-07 lb1 = -2.892018034e-13
+ keta = -1.746390476e-02 lketa = 8.039550078e-08 pketa = 1.110223025e-28
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -6.945600321e-01 lpclm = 5.993548011e-06 wpclm = 6.661338148e-22 ppclm = -1.776356839e-27
+ pdiblc1 = 0.39
+ pdiblc2 = -1.643357236e-03 lpdiblc2 = 2.567139102e-08 ppdiblc2 = -2.775557562e-29
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 6.390114615e+08 lpscbe1 = 2.870431763e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.862692334e-01 lkt1 = -3.884989683e-8
+ kt2 = -9.795153463e-03 lkt2 = -8.595216188e-8
+ at = 140000.0
+ ute = -1.231004634e+00 lute = -2.719492778e-7
+ ua1 = 1.515902718e-09 lua1 = -2.056269539e-15 wua1 = -3.308722450e-30
+ ub1 = -1.027457992e-18 lub1 = 1.411361252e-24
+ uc1 = -7.120287721e-11 luc1 = 4.117620565e-16 wuc1 = -5.169878828e-32 puc1 = 2.067951531e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 7.723053184e-04 ltvoff = -5.428361298e-09 ptvoff = 3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.147 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.326686961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.532798377e-8
+ k1 = 5.591506344e-01 lk1 = 2.756355115e-8
+ k2 = -3.874939645e-02 lk2 = -3.132893600e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.564204000e-01 ldsub = -1.178607824e-6
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.381492365e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.493671045e-8
+ nfactor = 2.371796068e+00 lnfactor = 3.545660917e-7
+ eta0 = 1.585514060e-01 leta0 = -3.123310732e-7
+ etab = -1.386707260e-01 letab = 2.730441458e-7
+ u0 = 3.007940389e-02 lu0 = -1.842556898e-9
+ ua = -7.055192805e-10 lua = 5.631706405e-16
+ ub = 1.674767488e-18 lub = -1.495653328e-24
+ uc = 3.557531560e-11 luc = 3.006628558e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.610603794e+00 la0 = -1.513332445e-6
+ ags = 3.267882410e-01 lags = 2.957519899e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.196129051e-08 lb0 = -9.782052066e-15
+ b1 = -1.129227465e-08 lb1 = 2.162313200e-13
+ keta = 5.179224004e-04 lketa = 8.897310460e-9
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.116334728e+00 lpclm = -1.206815837e-6
+ pdiblc1 = 0.39
+ pdiblc2 = 2.474187624e-03 lpdiblc2 = 9.299472665e-9
+ pdiblcb = -3.735085000e-02 lpdiblcb = 4.910865932e-8
+ drout = 0.56
+ pscbe1 = 6.234654264e+08 lpscbe1 = 3.488563261e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.587107910e-01 lkt1 = -1.484260119e-7
+ kt2 = -1.476078455e-02 lkt2 = -6.620813734e-8
+ at = 1.702645228e+05 lat = -1.203358588e-1
+ ute = -8.735426920e-01 lute = -1.693266573e-6
+ ua1 = 2.140334125e-09 lua1 = -4.539093737e-15
+ ub1 = -1.486104833e-18 lub1 = 3.235003467e-24 pub1 = -6.162975822e-45
+ uc1 = 8.417239227e-12 luc1 = 9.518164525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 4.235647164e-04 ltvoff = -4.041721236e-09 ptvoff = 3.469446952e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.148 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.382515671e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.429547149e-8
+ k1 = 5.915575913e-01 lk1 = -3.647700292e-8
+ k2 = -6.622449231e-02 lk2 = 2.296559004e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.26
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.732988774e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -5.321641882e-8
+ nfactor = 3.025795458e+00 lnfactor = -9.378256468e-07 wnfactor = 7.105427358e-21
+ eta0 = -1.482776250e-03 leta0 = 3.918235528e-09 peta0 = 3.469446952e-30
+ etab = 8.137340700e-02 letab = -1.617929870e-07 wetab = 2.775557562e-23 petab = -3.122502257e-29
+ u0 = 3.232676302e-02 lu0 = -6.283644175e-9
+ ua = 2.754445177e-10 lua = -1.375347236e-15
+ ub = 6.147365314e-20 lub = 1.692434697e-24
+ uc = 6.175884023e-11 luc = -2.167592006e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.666551942e+04 lvsat = 6.589387108e-3
+ a0 = 4.980764928e-01 la0 = 6.851728046e-7
+ ags = -2.786400028e-01 lags = 1.492160538e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -7.103458252e-08 lb0 = 1.542290805e-13 wb0 = -2.646977960e-29 pb0 = -2.646977960e-35
+ b1 = 1.871293712e-07 lb1 = -1.758768375e-13
+ keta = 7.110305558e-02 lketa = -1.305885123e-07 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.496432008e-01 lpclm = 7.034980908e-7
+ pdiblc1 = 4.247813265e-01 lpdiblc1 = -6.873263151e-8
+ pdiblc2 = 9.606198839e-03 lpdiblc2 = -4.794351448e-9
+ pdiblcb = -2.451476819e-02 lpdiblcb = 2.374281595e-8
+ drout = 2.088804448e-01 ldrout = 6.938599933e-7
+ pscbe1 = 8.645253716e+08 lpscbe1 = -1.275109097e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.328986640e-06 lalpha0 = 1.059008642e-11 walpha0 = 5.293955920e-28 palpha0 = -6.670384460e-33
+ alpha1 = 0.85
+ beta0 = 1.034200586e+01 lbeta0 = 6.952034876e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.915711146e-01 lkt1 = 1.141240567e-7
+ kt2 = -6.889893246e-02 lkt2 = 4.077620572e-8
+ at = 1.549379515e+05 lat = -9.004846934e-2
+ ute = -2.370540520e+00 lute = 1.265004727e-6
+ ua1 = -1.560482787e-09 lua1 = 2.774223792e-15 wua1 = -1.240770919e-30 pua1 = -1.654361225e-36
+ ub1 = 9.526220239e-19 lub1 = -1.584252469e-24 wub1 = 7.703719778e-40 pub1 = -3.851859889e-46
+ uc1 = 7.177850760e-11 luc1 = -3.002883819e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.016254171e-03 ltvoff = 7.796927017e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.149 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.489274262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.387438106e-8
+ k1 = 6.296133047e-01 lk1 = -7.362455483e-8
+ k2 = -7.127821251e-02 lk2 = 2.789870827e-08 pk2 = 5.551115123e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.120939287e-01 ldsub = 4.676284081e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.289427140e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.099533237e-9
+ nfactor = 2.132370221e+00 lnfactor = -6.572110951e-8
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = -2.636779683e-22 peta0 = -4.267419751e-28
+ etab = -1.641277800e-01 letab = 7.784955966e-8
+ u0 = 2.990485012e-02 lu0 = -3.919527800e-9
+ ua = -8.304373631e-10 lua = -2.958561202e-16
+ ub = 1.698955783e-18 lub = 9.402944032e-26
+ uc = 2.718870035e-11 luc = 1.206923800e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.039288954e+03 lvsat = 8.732052794e-2
+ a0 = 1.024210589e+00 la0 = 1.715943727e-7
+ ags = 2.291547500e+00 lags = -1.016692010e-6
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.697793345e-07 lb0 = -8.083805320e-14
+ b1 = 1.357375676e-08 lb1 = -6.462954249e-15
+ keta = -1.155907111e-01 lketa = 5.164999439e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.268894400e+00 lpclm = -3.890432980e-7
+ pdiblc1 = 6.603681753e-01 lpdiblc1 = -2.986974357e-7
+ pdiblc2 = 9.120988833e-03 lpdiblc2 = -4.320720495e-9
+ pdiblcb = 8.971602892e-02 lpdiblcb = -8.776197741e-08 wpdiblcb = -8.413408858e-23 ppdiblcb = 1.023486851e-28
+ drout = 8.432395256e-01 ldrout = 7.463925761e-8
+ pscbe1 = 1.016674454e+09 lpscbe1 = -2.760291061e+02 wpscbe1 = -1.907348633e-12
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.062680640e-06 lalpha0 = -1.505866109e-12
+ alpha1 = 0.85
+ beta0 = 1.693644131e+01 lbeta0 = 5.149690275e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.705693353e-01 lkt1 = -3.990136189e-9
+ kt2 = -1.799095058e-02 lkt2 = -8.916908084e-9
+ at = 1.122373800e+05 lat = -4.836690427e-02 wat = -2.328306437e-16
+ ute = -8.501885196e-01 lute = -2.190655934e-7
+ ua1 = 1.709985088e-09 lua1 = -4.181976374e-16 wua1 = 3.308722450e-30
+ ub1 = -7.070069558e-19 lub1 = 3.577112438e-26
+ uc1 = 7.460704526e-11 luc1 = -3.278987563e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.627520928e-04 ltvoff = -9.319638031e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.150 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.355705950e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -2.737955077e-8
+ k1 = 8.414013971e-02 lk1 = 1.860948561e-7
+ k2 = 1.046361009e-01 lk2 = -5.586042927e-08 wk2 = 1.110223025e-22 pk2 = -1.387778781e-29
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.761425679e-01 ldsub = 6.388057796e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-2.701903262e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 2.073900634e-8
+ nfactor = 8.725247214e-01 lnfactor = 5.341366871e-7
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.860778692e-02 letab = -1.868014223e-08 wetab = 2.775557562e-23 petab = 5.637851297e-30
+ u0 = 1.581860078e-02 lu0 = 2.787442612e-9
+ ua = -1.703807103e-09 lua = 1.199866543e-16
+ ub = 1.993090003e-18 lub = -4.601845039e-26
+ uc = 1.633443547e-11 luc = 1.723734426e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.620406891e+05 lvsat = 7.291599488e-3
+ a0 = 1.280215623e+00 la0 = 4.970115984e-8
+ ags = -8.330949999e-01 lags = 4.710627709e-07 wags = 4.440892099e-22 pags = 4.440892099e-28
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 6.166340672e-02 lketa = -3.274707227e-08 wketa = -2.775557562e-23 pketa = 2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.446949625e-01 lpclm = -9.183947451e-8
+ pdiblc1 = -2.599865133e-01 lpdiblc1 = 1.395165643e-07 wpdiblc1 = -1.110223025e-22 ppdiblc1 = 2.775557562e-29
+ pdiblc2 = -7.515255684e-03 lpdiblc2 = 3.600394425e-09 wpdiblc2 = 2.168404345e-25 ppdiblc2 = 3.794707604e-31
+ pdiblcb = -8.674421609e-02 lpdiblcb = -3.742902196e-9
+ drout = 1.449262700e+00 ldrout = -2.139101923e-7
+ pscbe1 = 1.163107023e+08 lpscbe1 = 1.526664890e+2
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 7.408183449e-06 lalpha0 = -1.670372435e-12
+ alpha1 = 0.85
+ beta0 = 2.136300371e+01 lbeta0 = -1.592676687e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.133121573e-01 lkt1 = 1.636126010e-8
+ kt2 = -4.380991832e-02 lkt2 = 3.376431938e-9
+ at = -5.685532692e+03 lat = 7.780439669e-3
+ ute = -1.302351205e+00 lute = -3.774660968e-9
+ ua1 = 1.605522255e-09 lua1 = -3.684591218e-16
+ ub1 = -1.843635241e-18 lub1 = 5.769607696e-25
+ uc1 = -1.222035414e-10 luc1 = 6.091872988e-17 wuc1 = -1.033975766e-31 puc1 = -3.231174268e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.228278134e-03 ltvoff = 9.561659042e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.151 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.703710179e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.263557920e-8
+ k1 = 9.070734896e-01 lk1 = 6.820322085e-17
+ k2 = -1.527159821e-01 lk2 = 2.336141377e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 4.586300001e-01 ldsub = -1.033750863e-17
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999996e-03 lcdscd = 7.217039466e-19
+ cit = 0.0
+ voff = {-1.136835598e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.465280779e-8
+ nfactor = 3.720571922e+00 lnfactor = -1.099093146e-7
+ eta0 = 2.242428860e-03 leta0 = -3.501238375e-10
+ etab = -4.399800002e-02 letab = 2.944755551e-18
+ u0 = 2.203500696e-02 lu0 = 1.381689384e-9
+ ua = -1.155463028e-09 lua = -4.013681436e-18
+ ub = 1.295395749e-18 lub = 1.117553374e-25
+ uc = 1.272578803e-10 luc = -7.846439865e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.854040931e+05 lvsat = 2.008292775e-3
+ a0 = 1.499999999e+00 la0 = 2.083488937e-16
+ ags = 1.250000000e+00 lags = 4.460964931e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -2.083869161e-01 lketa = 2.832102752e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.706266759e-01 lpclm = -2.986276845e-8
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566924534e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563599912e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889155499e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866149902e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 2.863680696e-09 lalpha0 = 4.236956351e-15
+ alpha1 = 0.85
+ beta0 = 1.533904646e+01 lbeta0 = -2.304430895e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.618011205e-01 lkt1 = 4.712760272e-9
+ kt2 = -2.887893901e-02 lkt2 = 1.131983396e-18
+ at = -2.704237011e+04 lat = 1.260998945e-2
+ ute = -1.326367013e+00 lute = 1.656177765e-9
+ ua1 = -2.384733737e-11 lua1 = 2.135940608e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034187072e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393363028e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.152 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 5.2e-07 wmax = 5.4e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {2.077259316e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 4.398637400e-08 wvth0 = 2.753432640e-07 pvth0 = -4.299099587e-14
+ k1 = 0.90707349
+ k2 = -1.907081280e-01 lk2 = 8.268083064e-09 wk2 = 1.937288518e-08 pk2 = -3.024804800e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.467965459e+00 ldsub = -3.137296012e-07 wdsub = -1.017279859e-06 pdsub = 1.588340081e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000001e-03 lcdscd = -1.335112576e-19
+ cit = 0.0
+ voff = {-2.075300001e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.749089762e-17
+ nfactor = 9.841048692e+00 lnfactor = -1.065536076e-06 wnfactor = -3.293789136e-06 pnfactor = 5.142790605e-13
+ eta0 = -1.136614629e-02 leta0 = 1.774664653e-09 weta0 = 4.276876273e-09 peta0 = -6.677743538e-16
+ etab = -0.043998
+ u0 = 1.847344735e-02 lu0 = 1.937777056e-09 wu0 = 3.205098134e-09 pu0 = -5.004312023e-16
+ ua = -1.477932599e-09 lua = 4.633542753e-17 wua = 1.398486904e-16 pua = -2.183541512e-23
+ ub = 6.883164335e-18 lub = -7.606964985e-25 wub = -2.980183442e-24 pub = 4.653139219e-31
+ uc = -2.014268208e-10 luc = 4.347307463e-17 wuc = 1.186133774e-16 puc = -1.851981829e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.068854253e+05 lvsat = -1.695931651e-02 wvsat = -3.771236119e-02 pvsat = 5.888257227e-9
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -8.229130756e-01 lketa = 1.242706840e-07 wketa = 4.029564638e-07 pketa = -6.291601043e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.088139166e-03 lpclm = 2.674254852e-08 wpclm = 1.207637111e-07 ppclm = -1.885556280e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.000000006e-08 lalpha0 = -9.450452472e-24 walpha0 = 2.191735868e-22 palpha0 = -3.422087222e-29
+ alpha1 = 0.85
+ beta0 = 1.391835560e+01 lbeta0 = -8.622102722e-09 wbeta0 = 3.967670636e-17 pbeta0 = -6.210143511e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.923331857e-01 lkt1 = -6.133685191e-09 wkt1 = -8.154366071e-17 pkt1 = 1.273181560e-23
+ kt2 = -0.028878939
+ at = 5.372048692e+04 lat = 1.022242941e-11 wat = -2.588424832e-11 pat = 4.041474313e-18
+ ute = -1.132927148e+00 lute = -2.854674899e-08 wute = -2.218108973e-07 pute = 3.463266627e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.0
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.153 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.154 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.700954295e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 7.609623444e-07 wvth0 = 1.049421690e-08 pvth0 = -2.096339040e-13
+ k1 = 8.217577412e-01 lk1 = -5.068944934e-06 wk1 = -9.974569897e-08 pk1 = 1.992533648e-12
+ k2 = -1.477861012e-01 lk2 = 2.122788586e-06 wk2 = 4.288599792e-08 pk2 = -8.566965270e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.763387208e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 5.931090735e-07 wvoff = 1.056299746e-08 pvoff = -2.110078738e-13
+ nfactor = 2.315264128e+00 lnfactor = 5.927036852e-06 wnfactor = 1.350000115e-07 pnfactor = -2.696778590e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 1.961436369e-02 lu0 = 1.041363222e-07 wu0 = 1.540117488e-09 pu0 = -3.076559639e-14
+ ua = -1.616986101e-09 lua = 1.124990859e-14 wua = 1.786897104e-16 pua = -3.569529956e-21
+ ub = 1.862903844e-18 lub = -5.317724193e-24 wub = -8.470113711e-26 pub = 1.692001434e-30
+ uc = 6.326296240e-11 luc = -2.941678276e-16 wuc = 2.025059733e-20 puc = -4.045286864e-25
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.060774878e+00 la0 = 6.029299683e-06 wa0 = 1.572399322e-07 pa0 = -3.141046271e-12
+ ags = 3.186892585e-01 lags = 5.231898148e-07 wags = 1.036354099e-09 pags = -2.070235042e-14
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 7.598262010e-08 lb0 = -1.504495294e-12 wb0 = -3.570742562e-14 pb0 = 7.132963903e-19
+ b1 = 1.199723230e-07 lb1 = -1.800835136e-12 wb1 = -5.868384865e-14 pb1 = 1.172276542e-18
+ keta = -5.263483841e-03 lketa = 1.432056911e-08 wketa = 1.239813041e-09 pketa = -2.476667393e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 5.695623324e-02 lpclm = -8.006681662e-07 wpclm = -3.175293662e-08 ppclm = 6.343009803e-13
+ pdiblc1 = 0.39
+ pdiblc2 = 3.210332764e-03 lpdiblc2 = -4.494641196e-08 wpdiblc2 = -1.266279500e-09 ppdiblc2 = 2.529537151e-14
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -1.041850928e+08 lpscbe1 = 6.575846183e+03 wpscbe1 = 1.432680922e+01 ppscbe1 = -2.861942893e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.009236635e-01 lkt1 = 2.905262004e-07 wkt1 = 8.433778183e-09 pkt1 = -1.684743000e-13
+ kt2 = -6.178975046e-02 lkt2 = 6.446662545e-07 wkt2 = 1.253822047e-08 pkt2 = -2.504651974e-13
+ at = 2.357796851e+05 lat = -1.214143255e+00 wat = -1.786817412e-02 pat = 3.569370762e-7
+ ute = -6.094748567e-01 lute = -1.010642947e-05 wute = -1.935718863e-07 pute = 3.866818326e-12
+ ua1 = 1.606117716e-09 lua1 = -9.690777475e-15 wua1 = -2.744551544e-16 pua1 = 5.482553491e-21
+ ub1 = -8.876086396e-19 lub1 = 6.355180732e-24 wub1 = 2.404937115e-25 pub1 = -4.804135088e-30
+ uc1 = 1.677082470e-10 luc1 = -2.674602552e-15 wuc1 = -4.686523553e-17 puc1 = 9.361863187e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.027033080e-04 ltvoff = -4.819308890e-09 wtvoff = -2.951822364e-11 ptvoff = 5.896600499e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.155 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.432776777e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(1))} lvth0 = 1.772507799e-07 wvth0 = -9.561110831e-09 pvth0 = -4.966988252e-14
+ k1 = -2.040130716e-01 lk1 = 3.112742574e-06 wk1 = 3.052782980e-07 pk1 = -1.237992835e-12
+ k2 = 2.830316823e-01 lk2 = -1.313472646e-06 wk2 = -1.289792910e-07 pk2 = 5.141243914e-13
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.443027856e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.375860969e-07 wvoff = -3.328537950e-09 pvoff = -1.002070981e-13
+ nfactor = 4.032210339e+00 lnfactor = -7.767559633e-06 wnfactor = -5.859982402e-07 pnfactor = 3.054001521e-12
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 3.225074892e-02 lu0 = 3.346795085e-09 wu0 = -2.974451048e-09 pu0 = 5.243216229e-15
+ ua = -1.865050936e-11 lua = -1.498633460e-15 wua = -4.563776808e-16 pua = 1.495853925e-21
+ ub = 9.153859060e-19 lub = 2.239807743e-24 wub = 3.393646320e-25 pub = -1.690404813e-30
+ uc = -7.681406779e-11 luc = 8.231056157e-16 wuc = 4.115715172e-17 puc = -3.285180466e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 2.175462013e+00 la0 = -2.861596503e-06 wa0 = -3.648315134e-07 pa0 = 1.023066581e-12
+ ags = 1.893441793e-01 lags = 1.554863758e-06 wags = 8.174241992e-08 pags = -6.644249075e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -3.580537256e-07 lb0 = 1.957437628e-12 wb0 = 1.661800130e-13 pb0 = -8.969852767e-19
+ b1 = -1.609955113e-07 lb1 = 4.402025214e-13 wb1 = 1.318443334e-13 pb1 = -3.474021506e-19
+ keta = -1.077482467e-02 lketa = 5.827977310e-08 wketa = -3.185888443e-09 pketa = 1.053332301e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.008746810e+00 lpclm = 1.567566024e-05 wpclm = 6.259235070e-07 ppclm = -4.611415778e-12
+ pdiblc1 = 0.39
+ pdiblc2 = -3.884875667e-03 lpdiblc2 = 1.164593544e-08 wpdiblc2 = 1.067594881e-09 ppdiblc2 = 6.680072035e-15
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 1.061386927e+09 lpscbe1 = -2.720914767e+03 wpscbe1 = -2.011698316e+02 ppscbe1 = 1.432636225e-3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.995756302e-01 lkt1 = 2.797741037e-07 wkt1 = 6.337597304e-09 pkt1 = -1.517548762e-13
+ kt2 = 2.322492653e-02 lkt2 = -3.342237117e-08 wkt2 = -1.572686974e-08 pkt2 = -2.501899378e-14
+ at = 2.745213476e+04 lat = 4.475056187e-01 wat = 5.360452235e-02 pat = -2.131388711e-7
+ ute = -2.827302572e+00 lute = 7.583266016e-06 wute = 7.602879747e-07 pute = -3.741297650e-12
+ ua1 = -1.784648604e-09 lua1 = 1.735443584e-14 wua1 = 1.571993185e-15 pua1 = -9.244969580e-21
+ ub1 = 1.459670687e-18 lub1 = -1.236703841e-23 wub1 = -1.184574622e-24 pub1 = 6.562403748e-30
+ uc1 = -2.939811106e-10 luc1 = 1.007894554e-15 wuc1 = 1.061052626e-16 puc1 = -2.839271782e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 2.303094330e-03 ltvoff = -1.838185894e-08 wtvoff = -7.290872521e-10 ptvoff = 6.169517762e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.156 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.633332245e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 9.750719844e-08 wvth0 = -1.460496290e-08 pvth0 = -2.961484072e-14
+ k1 = 6.989797175e-01 lk1 = -4.776795624e-07 wk1 = -6.659807534e-08 pk1 = 2.406382006e-13
+ k2 = -8.489741207e-02 lk2 = 1.494634718e-07 wk2 = 2.197946918e-08 pk2 = -8.610816957e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.971797010e+00 ldsub = -5.613496914e-06 wdsub = -5.312338023e-07 pdsub = 2.112257846e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-6.210270039e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -3.868662210e-07 wvoff = -8.384779633e-08 pvoff = 2.199484238e-13
+ nfactor = 9.180969716e-01 lnfactor = 4.614578636e-06 wnfactor = 6.923707129e-07 pnfactor = -2.028967295e-12
+ eta0 = 4.541262075e-01 leta0 = -1.487576682e-06 weta0 = -1.407769576e-07 peta0 = 5.597483292e-13
+ etab = -3.970663072e-01 letab = 1.300460118e-06 wetab = 1.230691642e-07 petab = -4.893397343e-13
+ u0 = 3.379753822e-02 lu0 = -2.803449534e-09 wu0 = -1.770880455e-09 pu0 = 4.576558666e-16
+ ua = -1.503415702e-09 lua = 4.404994874e-15 wua = 3.800237035e-16 pua = -1.829791730e-21
+ ub = 3.565806593e-18 lub = -8.298625364e-24 wub = -9.006678870e-25 pub = 3.240133127e-30
+ uc = 1.888221299e-10 luc = -2.331000331e-16 wuc = -7.298869923e-17 puc = 1.253413806e-22
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.328186982e+05 lvsat = -1.005241527e+00 wvsat = -1.204129952e-01 pvsat = 4.787784451e-7
+ a0 = 4.495430831e+00 la0 = -1.208610804e-05 wa0 = -1.373991191e-06 pa0 = 5.035622705e-12
+ ags = -9.049205322e-02 lags = 2.667530676e-06 wags = 1.987430931e-07 pags = -1.129635496e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 4.814907387e-08 lb0 = 3.423200541e-13 wb0 = -1.723558983e-14 pb0 = -1.676998953e-19
+ b1 = -3.395835565e-07 lb1 = 1.150292877e-12 wb1 = 1.563592283e-13 pb1 = -4.448767066e-19
+ keta = 5.073748949e-02 lketa = -1.863015537e-07 wketa = -2.391867585e-08 pketa = 9.296970541e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 8.147361128e+00 lpclm = -2.470640615e-05 wpclm = -3.348751316e-06 ppclm = 1.119243187e-11
+ pdiblc1 = 0.39
+ pdiblc2 = 1.418717630e-02 lpdiblc2 = -6.021100098e-08 wpdiblc2 = -5.578685672e-09 ppdiblc2 = 3.310658741e-14
+ pdiblcb = -8.382487540e-02 lpdiblcb = 2.338957048e-07 wpdiblcb = 2.213474176e-08 ppdiblcb = -8.801074358e-14
+ drout = 0.56
+ pscbe1 = -4.080239783e+07 lpscbe1 = 1.661539887e+03 wpscbe1 = 3.163788079e+02 ppscbe1 = -6.252075519e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -8.194415328e-02 lkt1 = -5.855582466e-07 wkt1 = -8.419076773e-08 pkt1 = 2.081982150e-13
+ kt2 = 1.434144464e-01 lkt2 = -5.113122478e-07 wkt2 = -7.533601533e-08 pkt2 = 2.119950759e-13
+ at = 2.841444747e+05 lat = -5.731380349e-01 wat = -5.423897122e-02 pat = 2.156615261e-7
+ ute = 1.909014365e+00 lute = -1.124897427e-05 wute = -1.325281840e-06 pute = 4.551211572e-12
+ ua1 = 1.141786848e-08 lua1 = -3.514056761e-14 wua1 = -4.418722615e-15 pua1 = 1.457493118e-20
+ ub1 = -7.308256149e-18 lub1 = 2.249543113e-23 wub1 = 2.772985873e-24 pub1 = -9.173395008e-30
+ uc1 = -1.786418358e-10 luc1 = 5.492899110e-16 wuc1 = 8.909287036e-17 puc1 = -2.162835930e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -4.156850401e-03 ltvoff = 7.303759866e-09 wtvoff = 2.181569273e-09 ptvoff = -5.403648430e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.157 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.078713948e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 9.493716740e-09 wvth0 = -3.315867078e-08 pvth0 = 7.049809357e-15
+ k1 = 4.780953274e-01 lk1 = -4.118196720e-08 wk1 = 5.404003399e-08 pk1 = 2.240889795e-15
+ k2 = -4.543748903e-02 lk2 = 7.148529733e-08 wk2 = -9.900475495e-09 pk2 = -2.310906322e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -1.970753219e+00 ldsub = 2.177518524e-06 wdsub = 1.062467605e-06 pdsub = -1.037112878e-12
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.085645523e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -9.743768276e-08 wvoff = 1.679640617e-08 pvoff = 2.106179203e-14
+ nfactor = 4.802023813e+00 lnfactor = -3.060589016e-06 wnfactor = -8.459855933e-07 pnfactor = 1.011033983e-12
+ eta0 = -5.926323793e-01 leta0 = 5.809606445e-07 weta0 = 2.815539152e-07 peta0 = -2.748349126e-13
+ etab = 9.069281548e-01 letab = -1.276410282e-06 wetab = -3.931968664e-07 petab = 5.308721543e-13
+ u0 = 3.149922292e-02 lu0 = 1.738334068e-09 wu0 = 3.941424525e-10 pu0 = -3.820723842e-15
+ ua = 2.205141162e-09 lua = -2.923617852e-15 wua = -9.190797770e-16 pua = 7.374134259e-22
+ ub = -3.228910931e-18 lub = 5.128660546e-24 wub = 1.567150951e-24 pub = -1.636612520e-30
+ uc = 1.124040642e-10 luc = -8.208754232e-17 wuc = -2.412140857e-17 puc = 2.877296827e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -8.890861700e+04 lvsat = -1.718509976e-01 wvsat = 7.885998084e-02 pvsat = 8.498794329e-8
+ a0 = -3.271981319e+00 la0 = 3.263354737e-06 wa0 = 1.795610675e-06 pa0 = -1.227941647e-12
+ ags = -2.579801431e+00 lags = 7.586744551e-06 wags = 1.096001767e-06 pags = -2.902740663e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -9.392010199e-07 lb0 = 2.293458119e-12 wb0 = 4.134920471e-13 pb0 = -1.018876285e-18
+ b1 = 4.956092053e-07 lb1 = -5.001616062e-13 wb1 = -1.469233923e-13 pb1 = 1.544509982e-19
+ keta = 2.707199972e-01 lketa = -6.210169064e-07 wketa = -9.507395617e-08 pketa = 2.335822164e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -8.849413375e+00 lpclm = 8.881531828e-06 wpclm = 4.286088664e-06 ppclm = -3.895050265e-12
+ pdiblc1 = 1.288078434e+00 lpdiblc1 = -1.774725125e-06 wpdiblc1 = -4.111728731e-07 ppdiblc1 = 8.125335167e-13
+ pdiblc2 = -3.255705279e-02 lpdiblc2 = 3.216195292e-08 wpdiblc2 = 2.008159781e-08 ppdiblc2 = -1.760162256e-14
+ pdiblcb = -2.268892823e-02 lpdiblcb = 1.130827587e-07 wpdiblcb = -8.696147089e-10 ppdiblcb = -4.255100660e-14
+ drout = -7.662332490e-01 ldrout = 2.620817268e-06 wdrout = 4.644291003e-07 pdrout = -9.177750646e-13
+ pscbe1 = 1.107322730e+09 lpscbe1 = -6.073115110e+02 wpscbe1 = -1.156400116e+02 ppscbe1 = 2.285203900e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -2.549388875e-05 lalpha0 = 5.043867542e-11 walpha0 = 9.604179906e-12 palpha0 = -1.897916566e-17
+ alpha1 = 0.85
+ beta0 = -2.895572869e+00 lbeta0 = 3.311129075e-05 wbeta0 = 6.304820470e-06 pbeta0 = -1.245918270e-11
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -5.576948819e-01 lkt1 = 3.545898952e-07 wkt1 = 7.912176010e-08 pkt1 = -1.145295505e-13
+ kt2 = -1.989770592e-01 lkt2 = 1.652999325e-07 wkt2 = 6.195387037e-08 pkt2 = -5.930840963e-14
+ at = 1.744165334e+05 lat = -3.563006999e-01 wat = -9.277297948e-03 pat = 1.268111449e-7
+ ute = -5.121844387e+00 lute = 2.644958824e-06 wute = 1.310396508e-06 pute = -6.572472969e-13
+ ua1 = -1.047559365e-08 lua1 = 8.123891057e-15 wua1 = 4.246106832e-15 pua1 = -2.547950225e-21
+ ub1 = 6.164193080e-18 lub1 = -4.127960800e-24 wub1 = -2.482177486e-24 pub1 = 1.211522491e-30
+ uc1 = 1.802776565e-10 luc1 = -1.599838187e-16 wuc1 = -5.167619164e-17 puc1 = 6.189521805e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -2.211137383e-03 ltvoff = 3.458766326e-09 wtvoff = 9.281936590e-11 ptvoff = -1.275994544e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.158 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.938860018e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.314536236e-08 wvth0 = -2.141296027e-08 pvth0 = -4.415601515e-15
+ k1 = 7.588584447e-01 lk1 = -3.152449535e-07 wk1 = -6.155713377e-08 pk1 = 1.150794467e-13
+ k2 = -7.581425847e-02 lk2 = 1.011371555e-07 wk2 = 2.160437041e-09 pk2 = -3.488215414e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.938772269e-01 ldsub = 6.454481925e-08 wdsub = 8.676287172e-09 pdsub = -8.469236255e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-3.571955599e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 4.764639450e-08 wvoff = 6.108452197e-08 pvoff = -2.216943217e-14
+ nfactor = 2.849888951e+00 lnfactor = -1.155039901e-06 wnfactor = -3.417412562e-07 pnfactor = 5.188229328e-13
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 4.336808690e-23 peta0 = -1.214306433e-29
+ etab = -7.805351919e-01 letab = 3.707834397e-07 wetab = 2.935837549e-07 petab = -1.395191343e-13
+ u0 = 5.261700169e-02 lu0 = -1.887549003e-08 wu0 = -1.081738898e-08 pu0 = 7.123255601e-15
+ ua = 8.824727399e-10 lua = -1.632513590e-15 wua = -8.158282496e-16 pua = 6.366258930e-22
+ ub = 9.981098225e-19 lub = 1.002513415e-24 wub = 3.338003158e-25 pub = -4.326945643e-31
+ uc = -1.672334365e-10 luc = 1.908766891e-16 wuc = 9.259976419e-17 puc = -8.516277042e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = -6.376868821e+05 lvsat = 3.638312230e-01 wvsat = 3.008423790e-01 pvsat = -1.316970669e-7
+ a0 = -7.660993235e-01 la0 = 8.172731101e-07 wa0 = 8.526923856e-07 pa0 = -3.075251604e-13
+ ags = 9.498328034e+00 lags = -4.203152431e-06 wags = -3.432459846e-06 pags = 1.517653742e-12
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.753340384e-06 lb0 = -1.310964477e-12 wb0 = -1.230503624e-12 pb0 = 5.858870735e-19
+ b1 = -3.275923799e-08 lb1 = 1.559785254e-14 wb1 = 2.206757140e-14 pb1 = -1.050716518e-20
+ keta = -6.875240046e-01 lketa = 3.143595604e-07 wketa = 2.724015329e-07 pketa = -1.251238375e-13
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 6.631978465e-01 lpclm = -4.040704387e-07 wpclm = 2.884823660e-07 ppclm = 7.157156668e-15
+ pdiblc1 = 6.058912244e-01 lpdiblc1 = -1.108817631e-06 wpdiblc1 = 2.594639114e-08 ppdiblc1 = 3.858456666e-13
+ pdiblc2 = 5.300944978e-03 lpdiblc2 = -4.792601592e-09 wpdiblc2 = 1.819418127e-09 ppdiblc2 = 2.247484731e-16
+ pdiblcb = 5.213717968e-01 lpdiblcb = -4.179945013e-07 wpdiblcb = -2.055898725e-07 ppdiblcb = 1.572838069e-13
+ drout = 2.793467272e+00 ldrout = -8.539345596e-07 wdrout = -9.288583713e-07 pdrout = 4.422629948e-13
+ pscbe1 = 1.831981422e+09 lpscbe1 = -1.314676947e+03 wpscbe1 = -3.883160333e+02 ppscbe1 = 4.946892711e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.556783204e-05 lalpha0 = -9.165868466e-12 walpha0 = -1.357649052e-11 palpha0 = 3.648321242e-18
+ alpha1 = 0.85
+ beta0 = 3.474735315e+01 lbeta0 = -3.633324486e-06 wbeta0 = -8.483016712e-06 pbeta0 = 1.975757531e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.102434031e-01 lkt1 = 1.542999846e-08 wkt1 = -2.873215566e-08 pkt1 = -9.249460571e-15
+ kt2 = -7.005837389e-02 lkt2 = 3.945776265e-08 wkt2 = 2.479877651e-08 pkt2 = -2.303998493e-14
+ at = -4.204198185e+05 lat = 2.243404773e-01 wat = 2.536950358e-01 pat = -1.298856171e-7
+ ute = -4.085857808e+00 lute = 1.633695028e-06 wute = 1.541091040e-06 pute = -8.824365344e-13
+ ua1 = -6.618614713e-09 lua1 = 4.358955067e-15 wua1 = 3.966762170e-15 pua1 = -2.275271845e-21
+ ub1 = 6.834047212e-18 lub1 = -4.781829534e-24 wub1 = -3.591668361e-24 pub1 = 2.294536477e-30
+ uc1 = 3.869173814e-10 luc1 = -3.616922933e-16 wuc1 = -1.487477915e-16 puc1 = 1.566503013e-22
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.405059855e-03 ltvoff = -3.975677982e-09 wtvoff = -2.699476810e-09 ptvoff = 1.449666276e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.159 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {7.582801055e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -5.512858863e-08 wvth0 = -5.844433107e-08 pvth0 = 1.321636725e-14
+ k1 = -6.361883992e-01 lk1 = 3.489870706e-07 wk1 = 3.430795172e-07 pk1 = -7.758262970e-14
+ k2 = 3.889507909e-01 lk2 = -1.201542160e-07 wk2 = -1.354139692e-07 pk2 = 3.062197333e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.125759715e-01 ldsub = 5.564167380e-08 wdsub = -1.735257434e-08 pdsub = 3.924041752e-15
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413313e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-3.282660694e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.387202260e-08 wvoff = 2.766043112e-08 pvoff = -6.255019251e-15
+ nfactor = -2.118204452e+00 lnfactor = 1.210448219e-06 wnfactor = 1.424430472e-06 pnfactor = -3.221150092e-13
+ eta0 = 9.325986798e-01 leta0 = -2.107371650e-7
+ etab = 3.636826934e-02 letab = -1.817370668e-08 wetab = 1.066641912e-09 petab = -2.412061354e-16
+ u0 = -7.489561147e-04 lu0 = 6.533963659e-09 wu0 = 7.890829134e-09 pu0 = -1.784400537e-15
+ ua = -3.788124322e-09 lua = 5.913258131e-16 wua = 9.927227740e-16 pua = -2.244903572e-22
+ ub = 4.292233931e-18 lub = -5.659376619e-25 wub = -1.095040869e-24 pub = 2.476281619e-31
+ uc = 3.612787256e-10 luc = -6.076697773e-17 wuc = -1.642907564e-16 puc = 3.715205449e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 6.508283590e+04 lvsat = 2.921726059e-02 wvsat = 4.617928026e-02 pvsat = -1.044279772e-8
+ a0 = 4.532065711e-01 la0 = 2.367176788e-07 wa0 = 3.938895252e-07 pa0 = -8.907260166e-14
+ ags = 1.466939411e-01 lags = 2.494972189e-07 wags = -4.666558364e-07 pags = 1.055276842e-13
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.322954847e-02 lketa = -2.405579330e-08 wketa = 1.830535488e-08 pketa = -4.139499730e-15
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -5.689893378e-01 lpclm = 1.826182384e-07 wpclm = 5.780559859e-07 ppclm = -1.307192684e-13
+ pdiblc1 = -3.604221043e+00 lpdiblc1 = 8.957683838e-07 wpdiblc1 = 1.592798710e-06 ppdiblc1 = -3.601891291e-13
+ pdiblc2 = -1.667822168e-02 lpdiblc2 = 5.672470903e-09 wpdiblc2 = 4.364155770e-09 ppdiblc2 = -9.868927293e-16
+ pdiblcb = -5.855669086e-01 lpdiblcb = 1.090588662e-07 wpdiblcb = 2.375802696e-07 ppdiblcb = -5.372545186e-14
+ drout = 1.449261983e+00 ldrout = -2.139100303e-07 wdrout = 3.413254115e-13 pdrout = -7.718596329e-20
+ pscbe1 = -2.485492668e+09 lpscbe1 = 7.410278960e+02 wpscbe1 = 1.239192113e+03 ppscbe1 = -2.802259477e-4
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.105748909e-05 lalpha0 = -7.018331815e-12 walpha0 = -1.126373859e-11 palpha0 = 2.547136789e-18
+ alpha1 = 0.85
+ beta0 = 3.869149493e+01 lbeta0 = -5.511272379e-06 wbeta0 = -8.253248456e-06 pbeta0 = 1.866356593e-12
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.207382264e-01 lkt1 = -2.718663834e-08 wkt1 = -9.171949695e-08 pkt1 = 2.074108016e-14
+ kt2 = 5.052406597e-02 lkt2 = -1.795587793e-08 wkt2 = -4.492957870e-08 pkt2 = 1.016019521e-14
+ at = 7.067492197e+04 lat = -9.487408107e-03 wat = -3.636911007e-02 pat = 8.224365075e-9
+ ute = -5.378324727e-02 lute = -2.861208247e-07 wute = -5.946704441e-07 pute = 1.344763955e-13
+ ua1 = 4.851948294e-09 lua1 = -1.102592921e-15 wua1 = -1.546214287e-15 pua1 = 3.496547140e-22
+ ub1 = -6.751768404e-18 lub1 = 1.686866370e-24 wub1 = 2.337655479e-24 pub1 = -5.286280594e-31
+ uc1 = -8.430044351e-10 luc1 = 2.239177608e-16 wuc1 = 3.433044912e-16 puc1 = -7.763350443e-23
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -5.608537609e-03 ltvoff = 1.268292261e-09 wtvoff = 6.573927431e-10 ptvoff = -1.486601653e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.25e-6
+ sbref = 1.24e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.160 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {2.319200945e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 6.390035881e-08 wvth0 = 1.611980827e-07 pvth0 = -3.645268963e-14
+ k1 = 9.070734896e-01 lk1 = 6.820277676e-17
+ k2 = -2.072877512e-01 lk2 = 1.467678295e-08 wk2 = 2.599155132e-08 pk2 = -5.877625449e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.844318224e+00 ldsub = -3.133539921e-07 wdsub = -6.599783585e-07 pdsub = 1.492448661e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999994e-03 lcdscd = 1.107712880e-18 wcdscd = 8.130007084e-19 pcdscd = -1.838485961e-25
+ cit = 0.0
+ voff = {-1.012324614e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.885622857e-07 wvoff = 4.280065586e-07 pvoff = -9.678769114e-14
+ nfactor = -4.823179794e+00 lnfactor = 1.822140524e-06 wnfactor = 4.069235155e-06 pnfactor = -9.202005610e-13
+ eta0 = 2.242427202e-03 leta0 = -3.501234117e-10 weta0 = 8.967860577e-16 peta0 = -2.027956119e-22
+ etab = -4.399800002e-02 letab = 2.944838817e-18
+ u0 = -3.174560466e-02 lu0 = 1.354342177e-08 wu0 = 2.561473726e-08 pu0 = -5.792414226e-15
+ ua = -1.020055485e-09 lua = -3.463420164e-17 wua = -6.449217553e-17 pua = 1.458400261e-23
+ ub = 6.725316299e-19 lub = 2.526073378e-25 wub = 2.966589683e-25 pub = -6.708527246e-32
+ uc = 2.485790391e-10 luc = -3.528152142e-17 wuc = -5.778308413e-17 puc = 1.306683551e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 7.550121294e+04 lvsat = 2.686129048e-02 wvsat = 5.234476356e-02 pvsat = -1.183703545e-8
+ a0 = 1.499999999e+00 la0 = 2.083475614e-16
+ ags = 1.250000000e+00 lags = 4.460964931e-17
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -5.556566672e-01 lketa = 1.068512200e-07 wketa = 1.653983316e-07 pketa = -3.740251712e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.856047518e-01 lpclm = -3.324985063e-08 wpclm = -7.133787964e-09 ppclm = 1.613206275e-15
+ pdiblc1 = 3.569721502e-01 lpdiblc1 = -3.566869022e-17
+ pdiblc2 = 8.406112094e-03 lpdiblc2 = 9.563565218e-19
+ pdiblcb = -1.032957700e-01 lpdiblcb = 2.831734847e-18
+ drout = 5.033266588e-01 ldrout = 1.889159940e-16
+ pscbe1 = 7.914198799e+08 lpscbe1 = 1.866316795e-8
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.841529940e-07 lalpha0 = -3.675908380e-14 walpha0 = -8.634483671e-14 palpha0 = 1.952567599e-20
+ alpha1 = 0.85
+ beta0 = 1.984497675e+01 lbeta0 = -1.249396142e-06 wbeta0 = -2.146093491e-06 pbeta0 = 4.853089976e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.723592454e-01 lkt1 = -1.551326758e-08 wkt1 = -4.259955513e-08 pkt1 = 9.633292999e-15
+ kt2 = -2.887893901e-02 lkt2 = 1.132025029e-18
+ at = -1.109726076e+05 lat = 3.158963765e-02 wat = 3.997446138e-02 pat = -9.039664800e-9
+ ute = -1.018204252e+00 lute = -6.803051626e-08 wute = -1.467723759e-07 pute = 3.319051800e-14
+ ua1 = -2.384733737e-11 lua1 = 2.135939962e-25
+ ub1 = 7.077531681e-19 lub1 = 3.034206331e-34
+ uc1 = 1.471862500e-10 luc1 = -4.393363028e-27
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.381383829e-03 ltvoff = 1.443060613e-09 wtvoff = 3.039338253e-09 ptvoff = -6.873037951e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.161 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 4.2e-07 wmax = 5.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {1.465520557e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -1.287090830e-07 wvth0 = -3.237216757e-07 pvth0 = 3.926074178e-14
+ k1 = 0.90707349
+ k2 = -1.042292523e-01 lk2 = -1.414358835e-09 wk2 = -2.181544669e-08 pk2 = 1.586767992e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -7.653070645e-01 ldsub = 9.410246186e-08 wdsub = 5.226696447e-07 pdsub = -3.540906255e-14
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.052000005e-03 lcdscd = -6.359062582e-19 wcdscd = -1.896999918e-18 pcdscd = 2.392799500e-25
+ cit = 0.0
+ voff = {4.998916816e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.754911788e-08 wvoff = -3.369322134e-07 pvoff = 2.264678897e-14
+ nfactor = 1.196065305e+01 lnfactor = -7.984200013e-07 wnfactor = -4.303318538e-06 pnfactor = 3.870564824e-13
+ eta0 = -1.136614502e-02 leta0 = 1.774664763e-09 weta0 = 4.276876208e-09 peta0 = -6.677744065e-16
+ etab = -0.043998
+ u0 = 1.424635325e-01 lu0 = -1.365689607e-08 wu0 = -5.584914762e-08 pu0 = 6.927030905e-15
+ ua = -1.793883530e-09 lua = 8.618821411e-17 wua = 2.903304318e-16 pua = -4.081658001e-23
+ ub = 8.336513898e-18 lub = -9.440161977e-25 wub = -3.672387679e-24 pub = 5.526257949e-31
+ uc = -4.845095256e-10 luc = 7.917999472e-17 wuc = 2.534405742e-16 puc = -3.552638160e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.461622170e+05 lvsat = -4.662583606e-02 wvsat = -1.516755901e-01 pvsat = 2.001788649e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.261698858e-02 lketa = 2.206317671e-08 wketa = 1.702702291e-08 pketa = -1.423641446e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.686070209e-02 lpclm = 3.115085549e-08 wpclm = 1.374092151e-07 ppclm = -2.095516005e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -3.930083952e-07 lalpha0 = 5.335658687e-14 walpha0 = 2.014712848e-13 palpha0 = -2.541278195e-20
+ alpha1 = 0.85
+ beta0 = 3.404518278e+00 lbeta0 = 1.317551282e-06 wbeta0 = 5.007551470e-06 pbeta0 = -6.316325119e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -4.010308949e-01 lkt1 = 2.019060909e-08 wkt1 = 9.939896227e-08 pkt1 = -1.253778751e-14
+ kt2 = -0.028878939
+ at = 2.495577075e+05 lat = -2.470212364e-02 wat = -9.327374313e-02 pat = 1.176517686e-8
+ ute = -1.851973592e+00 lute = 6.215089330e-08 wute = 1.206579809e-07 pute = -8.564988193e-15
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -6.955606043e-03 ltvoff = 1.532717373e-09 wtvoff = 3.312829958e-09 ptvoff = -7.300056959e-16
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.162 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.163 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.979846639e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.038432049e-7
+ k1 = 5.566754387e-01 lk1 = 2.263751931e-7
+ k2 = -3.381307583e-02 lk2 = -1.539520683e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.482666965e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.233849767e-8
+ nfactor = 2.674037632e+00 lnfactor = -1.239871451e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.370735110e-02 lu0 = 2.237424911e-8
+ ua = -1.142103671e-09 lua = 1.763592594e-15
+ ub = 1.637803688e-18 lub = -8.210928520e-25 wub = -1.540743956e-39
+ uc = 6.331678001e-11 luc = -2.952428955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.478652779e+00 la0 = -2.318286092e-6
+ ags = 3.214434537e-01 lags = 4.681716359e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.891276585e-08 lb0 = 3.911478418e-13 wb0 = -5.790264288e-30 pb0 = 9.926167351e-35
+ b1 = -3.598477475e-08 lb1 = 1.314585058e-12
+ keta = -1.968579909e-03 lketa = -5.149887994e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.742977677e-02 lpclm = 8.850382462e-7
+ pdiblc1 = 0.39
+ pdiblc2 = -1.549079328e-04 lpdiblc2 = 2.227809388e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.611043278e+07 lpscbe1 = 5.815261596e+03 ppscbe1 = -1.907348633e-18
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.785102125e-01 lkt1 = -1.572079458e-7
+ kt2 = -2.846841042e-02 lkt2 = -2.096536584e-8
+ at = 1.882935600e+05 lat = -2.655539625e-1
+ ute = -1.123907878e+00 lute = 1.699545360e-7
+ ua1 = 8.767308350e-10 lua1 = 4.879554061e-15
+ ub1 = -2.484770535e-19 lub1 = -6.412198755e-24
+ uc1 = 4.316007430e-11 luc1 = -1.866113153e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.242562293e-04 ltvoff = -3.252239379e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.164 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.178682486e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(1))} lvth0 = 4.524902983e-8
+ k1 = 6.072888189e-01 lk1 = -1.773240112e-7
+ k2 = -5.974126739e-02 lk2 = 5.285471378e-08 wk2 = -5.551115123e-23
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.531486457e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.127758856e-8
+ nfactor = 2.474872385e+00 lnfactor = 3.486976454e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.434590349e-02 lu0 = 1.728106839e-8
+ ua = -1.231511291e-09 lua = 2.476719931e-15
+ ub = 1.817275000e-18 lub = -2.252580446e-24
+ uc = 3.256440823e-11 luc = -4.995779590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205892612e+00 la0 = -1.427139067e-7
+ ags = 4.065813044e-01 lags = -2.108994399e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.358316642e-08 lb0 = -4.263736534e-13
+ b1 = 1.893915214e-07 lb1 = -4.830469315e-13
+ keta = -1.924158216e-02 lketa = 8.627293517e-08 pketa = 5.551115123e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.453042139e-01 lpclm = 3.420447988e-06 ppclm = 4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.047655494e-03 lpdiblc2 = 2.939876984e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.267617483e+08 lpscbe1 = 1.086432449e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.827329503e-01 lkt1 = -1.235268148e-7
+ kt2 = -1.857050812e-02 lkt2 = -9.991238073e-8
+ at = 1.699105100e+05 lat = -1.189282556e-1
+ ute = -8.067754816e-01 lute = -2.359536591e-6
+ ua1 = 2.393051059e-09 lua1 = -7.214822268e-15 pua1 = -6.617444900e-36
+ ub1 = -1.688432655e-18 lub1 = 5.073082956e-24
+ uc1 = -1.199775089e-11 luc1 = 2.533349999e-16 puc1 = -1.033975766e-37
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 3.654856960e-04 ltvoff = -1.985864012e-09 wtvoff = 2.168404345e-25
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.165 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.245193485e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.880335207e-8
+ k1 = 5.219899191e-01 lk1 = 1.618360153e-7
+ k2 = -2.648518619e-02 lk2 = -7.937598789e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.849350344e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.976645931e-7
+ nfactor = 2.758128419e+00 lnfactor = -7.775668681e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.909127947e-02 lu0 = -1.587191869e-9
+ ua = -4.934718209e-10 lua = -4.578253768e-16
+ ub = 1.172208475e-18 lub = 3.122917863e-25
+ uc = -5.151270940e-12 luc = 1.000048738e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.281137600e+04 lvsat = 2.671511067e-1
+ a0 = 8.439375600e-01 la0 = 1.296468606e-6
+ ags = 4.376838709e-01 lags = -3.345674742e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.344092944e-09 lb0 = -1.033560487e-13
+ b1 = 7.595380193e-08 lb1 = -3.200313110e-14
+ keta = -1.282833575e-02 lketa = 6.077299522e-08 wketa = 3.469446952e-24 pketa = -2.081668171e-29
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.522176873e-01 lpclm = 5.038391298e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -6.386343217e-04 lpdiblc2 = 2.777244603e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.056879617e-01 lkt1 = -3.225456744e-8
+ kt2 = -5.679713785e-02 lkt2 = 5.208189791e-8
+ at = 140000.0
+ ute = -1.613029847e+00 lute = 8.462404173e-7
+ ua1 = -3.252460382e-10 lua1 = 3.593496680e-15
+ ub1 = 6.117920260e-20 lub1 = -1.883611737e-24
+ uc1 = 5.812970886e-11 luc1 = -2.550131747e-17 wuc1 = -5.169878828e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.640847264e-03 ltvoff = -7.056875057e-09 ptvoff = 8.673617380e-31
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.166 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.197495320e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.822915813e-8
+ k1 = 6.217111102e-01 lk1 = -3.522662043e-8
+ k2 = -7.174880739e-02 lk2 = 1.007108346e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.639267377e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.146425849e-8
+ nfactor = 2.553748335e+00 lnfactor = -3.736840271e-7
+ eta0 = 1.556200357e-01 leta0 = -1.494354750e-7
+ etab = -1.380244775e-01 letab = 1.344256189e-7
+ u0 = 3.254668853e-02 lu0 = -8.415550098e-9
+ ua = -2.373880505e-10 lua = -9.638817346e-16
+ ub = 9.359201014e-19 lub = 7.792297471e-25
+ uc = 4.829946030e-11 luc = -5.621040407e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.206681920e+05 lvsat = 5.401136973e-2
+ a0 = 1.5
+ ags = 3.329123510e-01 lags = -1.275247019e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.596877049e-07 lb0 = -4.142884246e-13
+ b1 = 1.051483479e-07 lb1 = -8.969552433e-14
+ keta = 1.805323083e-02 lketa = -2.531802246e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.541215632e+00 lpclm = -1.469880848e-6
+ pdiblc1 = 1.953531031e-01 lpdiblc1 = 3.846487403e-7
+ pdiblc2 = 2.081142567e-02 lpdiblc2 = -1.461578972e-8
+ pdiblcb = -0.025
+ drout = 4.680248349e-01 ldrout = 1.817554350e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.474223732e-01 lkt1 = 5.021830556e-8
+ kt2 = -3.432961298e-02 lkt2 = 7.683013180e-9
+ at = 1.497613600e+05 lat = -1.928977490e-2
+ ute = -1.639359155e+00 lute = 8.982707095e-7
+ ua1 = 8.087803889e-10 lua1 = 1.352506233e-15
+ ub1 = -4.323953449e-19 lub1 = -9.082413048e-25
+ uc1 = 4.294397687e-11 luc1 = 4.507754196e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.964462374e-03 ltvoff = 6.770710992e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.167 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.369793193e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.141054242e-8
+ k1 = 5.952653582e-01 lk1 = -9.411969933e-9
+ k2 = -7.007272143e-02 lk2 = 8.434995606e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.169351653e-01 ldsub = 4.203713551e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.948584777e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.127067349e-8
+ nfactor = 1.941683786e+00 lnfactor = 2.237742136e-7
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = -1.630640067e-22 peta0 = 5.898059818e-29
+ etab = -0.0003125
+ u0 = 2.386891122e-02 lu0 = 5.514072691e-11
+ ua = -1.285657146e-09 lua = 5.937146704e-17
+ ub = 1.885211294e-18 lub = -1.474075602e-25
+ uc = 7.885796353e-11 luc = -3.545029551e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.618261931e+05 lvsat = 1.383556317e-2
+ a0 = 1.5
+ ags = 3.762869949e-01 lags = -1.698642534e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.168230143e-07 lb0 = 2.460780427e-13
+ b1 = 2.588712672e-08 lb1 = -1.232579297e-14
+ keta = 3.640521038e-02 lketa = -1.816720814e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.429863183e+00 lpclm = -3.850497131e-7
+ pdiblc1 = 6.748458678e-01 lpdiblc1 = -8.340140914e-8
+ pdiblc2 = 1.013619654e-02 lpdiblc2 = -4.195314257e-9
+ pdiblcb = -0.025
+ drout = 3.249506503e-01 ldrout = 3.214152972e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.127950400e-07 lalpha0 = 5.298417792e-13 walpha0 = 1.588186776e-28 palpha0 = -1.588186776e-34
+ alpha1 = 0.85
+ beta0 = 1.220304672e+01 lbeta0 = 1.617411747e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.866014421e-01 lkt1 = -9.151194823e-9
+ kt2 = -4.153609621e-03 lkt2 = -2.177287003e-8
+ at = 2.537953600e+05 lat = -1.208411075e-1
+ ute = 9.716893932e-03 lute = -7.114517882e-7
+ ua1 = 3.923378182e-09 lua1 = -1.687764798e-15
+ ub1 = -2.711103396e-18 lub1 = 1.316087658e-24
+ uc1 = -8.391965094e-12 luc1 = 5.461861525e-17 puc1 = -2.584939414e-38
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.769019187e-03 ltvoff = -1.230720203e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.168 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-7.962539828e-02+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.049982462e-07 wvth0 = 2.568444277e-07 pvth0 = -1.222928784e-13
+ k1 = 2.755733053e-01 lk1 = 1.428049254e-07 wk1 = -5.312266183e-16 pk1 = 2.529363385e-22
+ k2 = 9.547334747e-03 lk2 = -2.947497946e-08 wk2 = 7.348722109e-09 pk2 = -3.498991150e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.890254365e+00 ldsub = -7.546903751e-07 wdsub = -6.486327557e-07 pdsub = 3.088374058e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413326e-03 lcdscd = -1.441936607e-09 wcdscd = -4.822274524e-18 pcdscd = 2.296059176e-24
+ cit = 0.0
+ voff = {-1.675972920e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 6.939412324e-07 wvoff = 5.347782601e-07 pvoff = -2.546271817e-13
+ nfactor = -1.123616795e+01 lnfactor = 6.498223828e-06 wnfactor = 4.855356013e-06 pnfactor = -2.311809791e-12
+ eta0 = 9.253513184e-01 leta0 = -2.072863913e-07 weta0 = 2.727086470e-09 peta0 = -1.298464043e-15
+ etab = 3.920295698e-02 letab = -1.881473162e-08 wetab = -2.293703942e-17 petab = 1.092114778e-23
+ u0 = -1.808091525e-02 lu0 = 2.002896330e-08 wu0 = 1.441253338e-08 pu0 = -6.862325993e-15
+ ua = -1.064517984e-09 lua = -4.592084904e-17 wua = -3.212126641e-17 pua = 1.529409130e-23
+ ub = 2.920531487e-18 lub = -6.403607759e-25 wub = -5.788939296e-25 pub = 2.756322401e-31
+ uc = -8.683275570e-11 luc = 4.344102078e-17 wuc = 4.325528016e-18 puc = -2.059539608e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 9.266001192e+04 lvsat = 4.676807202e-02 wvsat = 3.580248531e-02 pvsat = -1.704685215e-8
+ a0 = 1.500000005e+00 la0 = -2.231342222e-15 wa0 = -1.622799672e-15 pa0 = 7.726734808e-22
+ ags = -1.093481874e+00 lags = 5.299456168e-07 wags = -3.474567301e-16 pags = 1.654362758e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 2.261106420e-01 lketa = -1.084927935e-07 wketa = -5.803514877e-08 pketa = 2.763262359e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 3.677243673e-01 lpclm = 1.206728138e-07 wpclm = 2.255874795e-07 ppclm = -1.074103202e-13
+ pdiblc1 = 6.287709947e-01 lpdiblc1 = -6.146350335e-08 wpdiblc1 = 2.778195451e-16 ppdiblc1 = -1.322800758e-22
+ pdiblc2 = -5.080122972e-03 lpdiblc2 = 3.049723249e-09 wpdiblc2 = -7.448985873e-18 ppdiblc2 = 3.546732786e-24
+ pdiblcb = 4.582196904e-02 lpdiblcb = -3.372088905e-08 wpdiblcb = -2.205591265e-17 ppdiblcb = 1.050159959e-23
+ drout = 1.449262894e+00 ldrout = -2.139102373e-07 wdrout = -1.471450517e-15 pdrout = 7.006102365e-22
+ pscbe1 = 8.077610965e+08 lpscbe1 = -3.695337436e+00 wpscbe1 = -1.453666687e-07 ppscbe1 = 6.921434402e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.436415553e-06 lalpha0 = -3.982475555e-13 walpha0 = -1.178617961e-13 palpha0 = 5.611824414e-20
+ alpha1 = 0.85
+ beta0 = 1.759308914e+01 lbeta0 = -9.489814890e-07 wbeta0 = -3.142981258e-07 pbeta0 = 1.496486524e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.556720410e-01 lkt1 = -7.149139618e-08 wkt1 = -7.857453133e-08 pkt1 = 3.741216305e-14
+ kt2 = -6.887994138e-02 lkt2 = 9.045666669e-09 wkt2 = -8.817280239e-18 pkt2 = 4.198211223e-24
+ at = 1.306347085e+05 lat = -6.219988757e-02 wat = -5.893089846e-02 pat = 2.805912227e-8
+ ute = -1.216531881e+00 lute = -1.275906013e-07 wute = -1.571490625e-07 pute = 7.482432602e-14
+ ua1 = 7.427581515e-10 lua1 = -1.733570997e-16 wua1 = -1.663665766e-24 pua1 = 7.921313156e-31
+ ub1 = -5.392589525e-19 lub1 = 2.819943316e-25 wub1 = -2.363318072e-33 pub1 = 1.125260585e-39
+ uc1 = 6.935515480e-11 luc1 = 1.760041257e-17 wuc1 = 3.421922117e-26 puc1 = -1.629297653e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.179989579e-02 ltvoff = 4.652989441e-09 wtvoff = 2.987089381e-09 ptvoff = -1.422260790e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.169 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {3.098120471e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -4.136044937e-07 wvth0 = -9.173015275e-07 pvth0 = 1.432237913e-13
+ k1 = 9.070734845e-01 lk1 = 8.554508213e-16 wk1 = 1.897239699e-15 pk1 = -2.962274870e-22
+ k2 = -6.846371117e-02 lk2 = -1.183387358e-08 wk2 = -2.624543611e-08 pk2 = 4.097857412e-15
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = -6.066036018e+00 ldsub = 1.044513307e-06 wdsub = 2.316545556e-06 pdsub = -3.616961569e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 2.051999950e-03 lcdscd = 7.765460150e-18 wcdscd = 1.722241447e-17 pcdscd = -2.689038228e-24
+ cit = 0.0
+ voff = {5.200911512e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -8.611699055e-07 wvoff = -1.909922358e-06 pvoff = 2.982076372e-13
+ nfactor = 5.207508359e+01 lnfactor = -7.818729352e-06 wnfactor = -1.734055719e-05 pnfactor = 2.707485237e-12
+ eta0 = 2.812619630e-02 leta0 = -4.391511347e-09 weta0 = -9.739594534e-09 peta0 = 1.520701332e-15
+ etab = -4.399800024e-02 letab = 3.693628736e-17 wetab = 8.191813894e-17 petab = -1.279036599e-23
+ u0 = 1.731222093e-01 lu0 = -2.320894646e-08 wu0 = -5.147333350e-08 pu0 = 8.036840399e-15
+ ua = -1.496323242e-09 lua = 5.172586476e-17 wua = 1.147188086e-16 pua = -1.791173590e-23
+ ub = -4.033564733e-18 lub = 9.322107271e-25 wub = 2.067478320e-24 pub = -3.228077950e-31
+ uc = 1.360709473e-10 luc = -6.965531008e-18 wuc = -1.544831434e-17 puc = 2.412038008e-24
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 5.544260154e+05 lvsat = -5.765384495e-02 wvsat = -1.278660190e-01 pvsat = 1.996448874e-8
+ a0 = 1.499999983e+00 la0 = 2.613244732e-15 wa0 = 5.795715907e-15 pa0 = -9.049196947e-22
+ ags = 1.249999996e+00 lags = 5.595195418e-16 wags = 1.240916703e-15 pags = -1.937512373e-22
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -6.669297466e-01 lketa = 9.345578777e-08 wketa = 2.072683885e-07 pketa = -3.236205710e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.507778499e+00 lpclm = -3.632704673e-07 wpclm = -8.056695698e-07 ppclm = 1.257940240e-13
+ pdiblc1 = 3.569721529e-01 lpdiblc1 = -4.473816873e-16 wpdiblc1 = -9.922134225e-16 ppdiblc1 = 1.549202988e-22
+ pdiblc2 = 8.406112023e-03 lpdiblc2 = 1.199532834e-17 wpdiblc2 = 2.660351106e-17 ppdiblc2 = -4.153767608e-24
+ pdiblcb = -1.032957702e-01 lpdiblcb = 3.551725580e-17 wpdiblcb = 7.877121178e-17 ppdiblcb = -1.229899516e-23
+ drout = 5.033266448e-01 ldrout = 2.369521024e-15 wdrout = 5.255178515e-15 pdrout = -8.205225388e-22
+ pscbe1 = 7.914198785e+08 lpscbe1 = 2.340879440e-07 wpscbe1 = 5.191669464e-07 ppscbe1 = -8.106064796e-14
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -1.163984368e-06 lalpha0 = 1.897964808e-13 walpha0 = 4.209349860e-13 palpha0 = -6.572310497e-20
+ alpha1 = 0.85
+ beta0 = 1.115844166e+01 lbeta0 = 5.061239535e-07 wbeta0 = 1.122493306e-06 pbeta0 = -1.752616149e-13
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.031350325e+00 lkt1 = 1.265309882e-07 wkt1 = 2.806233262e-07 pkt1 = -4.381540366e-14
+ kt2 = -2.887893909e-02 lkt2 = 1.419867002e-17 wkt2 = 3.149014383e-17 pkt2 = -4.916747565e-24
+ at = -5.640717012e+05 lat = 9.489824110e-02 wat = 2.104674945e-01 pat = -3.286155272e-8
+ ute = -2.899822368e+00 lute = 2.530619761e-07 wute = 5.612466518e-07 pute = -8.763080722e-14
+ ua1 = -2.384735316e-11 lua1 = 2.679052638e-24 wua1 = 5.941664344e-24 pua1 = -9.277077044e-31
+ ub1 = 7.077531456e-19 lub1 = 3.805723081e-33 wub1 = 8.440420337e-33 pub1 = -1.317853387e-39
+ uc1 = 1.471862504e-10 luc1 = -5.510429087e-26 wuc1 = -1.222117996e-25 puc1 = 1.908160917e-32
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 3.004745044e-02 ltvoff = -4.810202045e-09 wtvoff = -1.066817636e-08 ptvoff = 1.665686385e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.170 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.9e-07 wmax = 4.2e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-1.845492211e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 3.582714160e-07 wvth0 = 9.221528304e-07 pvth0 = -1.439812543e-13
+ k1 = 0.90707349
+ k2 = -1.469863474e+00 lk2 = 2.069750797e-07 wk2 = 4.920481293e-07 pk2 = -7.682642672e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.327233918e+00 ldsub = -4.221142877e-07 wdsub = -1.017279861e-06 pdsub = 1.588340084e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {3.866578765e+00+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -6.528325277e-07 wvoff = -1.603755963e-06 pvoff = 2.504040410e-13
+ nfactor = 3.541633038e+01 lnfactor = -5.217698260e-06 wnfactor = -1.312926772e-05 pnfactor = 2.049951344e-12
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 5.002217776e-01 lu0 = -7.428096467e-08 wu0 = -1.904671356e-07 pu0 = 2.973877668e-14
+ ua = -1.393966080e-09 lua = 3.574422705e-17 wua = 1.398486939e-16 pua = -2.183541567e-23
+ ub = 6.496925019e-18 lub = -7.119778210e-25 wub = -2.980183497e-24 pub = 4.653139304e-31
+ uc = -1.261952878e-10 luc = 3.398366988e-17 wuc = 1.186133762e-16 puc = -1.851981810e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 4.815522429e+05 lvsat = -4.627562560e-02 wvsat = -1.273640198e-01 pvsat = 1.988610860e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.038255850e+00 lketa = 1.514331602e-07 wketa = 4.029564649e-07 pketa = -6.291601060e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.737606982e-02 lpclm = 2.557100636e-08 wpclm = 1.207637141e-07 ppclm = -1.885556327e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.424179121e-07 lalpha0 = -1.417994553e-14 walpha0 = 2.955654554e-21 palpha0 = -4.614840902e-28
+ alpha1 = 0.85
+ beta0 = 1.671249328e+01 lbeta0 = -3.610634506e-07 wbeta0 = 2.044754410e-14 pbeta0 = -3.192596409e-21
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.368700706e-01 lkt1 = -1.312958075e-08 wkt1 = -1.018287676e-15 pkt1 = 1.589913756e-22
+ kt2 = -0.028878939
+ at = 1.675154536e+03 lat = 6.564790030e-03 wat = -3.270385787e-10 pat = 5.106249591e-17
+ ute = -9.418347041e-01 lute = -5.265038572e-08 wute = -2.218109000e-07 pute = 3.463266668e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 6.886122803e-02 ltvoff = -1.087043002e-08 wtvoff = -2.521568000e-08 ptvoff = 3.937075413e-15
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.171 nmos
* Model Flag Parameters
+ lmin = 2.0e-05 lmax = 0.0001 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.508189+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.56800772
+ k2 = -0.041519875
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-0.24664784+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 2.61197
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 0.0248274
+ ua = -1.0538187e-9
+ ub = 1.5967e-18
+ uc = 4.8537e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.3626
+ ags = 0.34488
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 6.6799e-10
+ b1 = 2.9823e-8
+ keta = -0.0045466
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.016875
+ pdiblc1 = 0.39
+ pdiblc2 = 0.00096032746
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 225000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.28638
+ kt2 = -0.029517931
+ at = 175000.0
+ ute = -1.1154
+ ua1 = 1.121e-9
+ ub1 = -5.6947e-19
+ uc1 = 3.3818362e-11
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 0.00036145
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.172 nmos
* Model Flag Parameters
+ lmin = 8.0e-06 lmax = 2.0e-05 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {4.979846639e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.038432049e-7
+ k1 = 5.566754387e-01 lk1 = 2.263751931e-7
+ k2 = -3.381307583e-02 lk2 = -1.539520683e-7
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.482666965e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 3.233849767e-8
+ nfactor = 2.674037632e+00 lnfactor = -1.239871451e-6
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.370735110e-02 lu0 = 2.237424911e-8
+ ua = -1.142103671e-09 lua = 1.763592594e-15 wua = 8.271806126e-31
+ ub = 1.637803688e-18 lub = -8.210928520e-25
+ uc = 6.331678001e-11 luc = -2.952428955e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.478652779e+00 la0 = -2.318286092e-6
+ ags = 3.214434537e-01 lags = 4.681716359e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -1.891276585e-08 lb0 = 3.911478418e-13 pb0 = 2.646977960e-35
+ b1 = -3.598477475e-08 lb1 = 1.314585058e-12 pb1 = 4.235164736e-34
+ keta = -1.968579909e-03 lketa = -5.149887994e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -2.742977677e-02 lpclm = 8.850382462e-07 ppclm = 1.110223025e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.549079328e-04 lpdiblc2 = 2.227809388e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = -6.611043278e+07 lpscbe1 = 5.815261596e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.785102125e-01 lkt1 = -1.572079458e-07 wkt1 = -2.220446049e-22
+ kt2 = -2.846841042e-02 lkt2 = -2.096536584e-8
+ at = 1.882935600e+05 lat = -2.655539625e-1
+ ute = -1.123907878e+00 lute = 1.699545360e-7
+ ua1 = 8.767308350e-10 lua1 = 4.879554061e-15
+ ub1 = -2.484770535e-19 lub1 = -6.412198755e-24
+ uc1 = 4.316007430e-11 luc1 = -1.866113153e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 5.242562293e-04 ltvoff = -3.252239379e-9
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.173 nmos
* Model Flag Parameters
+ lmin = 4.0e-06 lmax = 8.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.178682486e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope1/sqrt(1))} lvth0 = 4.524902983e-8
+ k1 = 6.072888189e-01 lk1 = -1.773240112e-7
+ k2 = -5.974126739e-02 lk2 = 5.285471378e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.531486457e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.127758856e-8
+ nfactor = 2.474872385e+00 lnfactor = 3.486976454e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.434590349e-02 lu0 = 1.728106839e-8
+ ua = -1.231511291e-09 lua = 2.476719931e-15
+ ub = 1.817275000e-18 lub = -2.252580446e-24
+ uc = 3.256440823e-11 luc = -4.995779590e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 80000.0
+ a0 = 1.205892612e+00 la0 = -1.427139067e-7
+ ags = 4.065813044e-01 lags = -2.108994399e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 8.358316642e-08 lb0 = -4.263736534e-13 pb0 = -1.058791184e-34
+ b1 = 1.893915215e-07 lb1 = -4.830469315e-13
+ keta = -1.924158216e-02 lketa = 8.627293517e-8
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -3.453042139e-01 lpclm = 3.420447988e-06 wpclm = 1.110223025e-22 ppclm = -4.440892099e-28
+ pdiblc1 = 0.39
+ pdiblc2 = -1.047655494e-03 lpdiblc2 = 2.939876984e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 5.267617483e+08 lpscbe1 = 1.086432449e+3
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.827329503e-01 lkt1 = -1.235268148e-7
+ kt2 = -1.857050812e-02 lkt2 = -9.991238073e-8
+ at = 1.699105100e+05 lat = -1.189282556e-1
+ ute = -8.067754816e-01 lute = -2.359536591e-6
+ ua1 = 2.393051059e-09 lua1 = -7.214822268e-15 wua1 = 1.654361225e-30
+ ub1 = -1.688432655e-18 lub1 = 5.073082956e-24
+ uc1 = -1.199775089e-11 luc1 = 2.533349999e-16
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 3.654856960e-04 ltvoff = -1.985864012e-09 wtvoff = 1.084202172e-25 ptvoff = 4.336808690e-31
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.174 nmos
* Model Flag Parameters
+ lmin = 2.0e-06 lmax = 4.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.245193485e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.880335207e-8
+ k1 = 5.219899191e-01 lk1 = 1.618360153e-7
+ k2 = -2.648518619e-02 lk2 = -7.937598789e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.56
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-2.849350344e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 1.976645931e-7
+ nfactor = 2.758128419e+00 lnfactor = -7.775668681e-7
+ eta0 = 0.08
+ etab = -0.07
+ u0 = 2.909127947e-02 lu0 = -1.587191869e-9
+ ua = -4.934718209e-10 lua = -4.578253768e-16
+ ub = 1.172208475e-18 lub = 3.122917863e-25
+ uc = -5.151270940e-12 luc = 1.000048738e-16
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.281137600e+04 lvsat = 2.671511067e-1
+ a0 = 8.439375600e-01 la0 = 1.296468606e-6
+ ags = 4.376838709e-01 lags = -3.345674742e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 2.344092944e-09 lb0 = -1.033560487e-13
+ b1 = 7.595380193e-08 lb1 = -3.200313110e-14
+ keta = -1.282833575e-02 lketa = 6.077299522e-08 wketa = 3.469446952e-24
+ dwg = 0.0
+ dwb = 0.0
+ pclm = -7.522176873e-01 lpclm = 5.038391298e-6
+ pdiblc1 = 0.39
+ pdiblc2 = -6.386343217e-04 lpdiblc2 = 2.777244603e-8
+ pdiblcb = -0.025
+ drout = 0.56
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.056879617e-01 lkt1 = -3.225456744e-8
+ kt2 = -5.679713785e-02 lkt2 = 5.208189791e-8
+ at = 140000.0
+ ute = -1.613029847e+00 lute = 8.462404173e-7
+ ua1 = -3.252460382e-10 lua1 = 3.593496680e-15
+ ub1 = 6.117920260e-20 lub1 = -1.883611737e-24
+ uc1 = 5.812970886e-11 luc1 = -2.550131747e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = 1.640847264e-03 ltvoff = -7.056875057e-09 wtvoff = -1.084202172e-25 ptvoff = 1.734723476e-30
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.175 nmos
* Model Flag Parameters
+ lmin = 1.0e-06 lmax = 2.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-09*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.197495320e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 2.822915813e-8
+ k1 = 6.217111102e-01 lk1 = -3.522662043e-8
+ k2 = -7.174880739e-02 lk2 = 1.007108346e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 8.528408000e-01 ldsub = -5.786932471e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.639267377e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.146425849e-8
+ nfactor = 2.553748335e+00 lnfactor = -3.736840271e-7
+ eta0 = 1.556200358e-01 leta0 = -1.494354750e-7
+ etab = -1.380244775e-01 letab = 1.344256189e-7
+ u0 = 3.254668853e-02 lu0 = -8.415550098e-9
+ ua = -2.373880505e-10 lua = -9.638817346e-16
+ ub = 9.359201014e-19 lub = 7.792297471e-25
+ uc = 4.829946030e-11 luc = -5.621040407e-18
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.206681920e+05 lvsat = 5.401136973e-2
+ a0 = 1.5
+ ags = 3.329123510e-01 lags = -1.275247019e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 1.596877049e-07 lb0 = -4.142884246e-13 wb0 = 5.293955920e-29 pb0 = 1.058791184e-34
+ b1 = 1.051483479e-07 lb1 = -8.969552433e-14
+ keta = 1.805323083e-02 lketa = -2.531802246e-10
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 2.541215632e+00 lpclm = -1.469880848e-6
+ pdiblc1 = 1.953531031e-01 lpdiblc1 = 3.846487403e-7
+ pdiblc2 = 2.081142567e-02 lpdiblc2 = -1.461578972e-8
+ pdiblcb = -0.025
+ drout = 4.680248349e-01 ldrout = 1.817554350e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 3.0e-8
+ alpha1 = 0.85
+ beta0 = 13.86
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.474223732e-01 lkt1 = 5.021830556e-8
+ kt2 = -3.432961298e-02 lkt2 = 7.683013180e-9
+ at = 1.497613600e+05 lat = -1.928977490e-2
+ ute = -1.639359155e+00 lute = 8.982707095e-7
+ ua1 = 8.087803889e-10 lua1 = 1.352506233e-15
+ ub1 = -4.323953449e-19 lub1 = -9.082413048e-25
+ uc1 = 4.294397687e-11 luc1 = 4.507754196e-18
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.964462374e-03 ltvoff = 6.770710992e-11
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 2.75e-6
+ sbref = 2.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.176 nmos
* Model Flag Parameters
+ lmin = 5.0e-07 lmax = 1.0e-06 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {5.369793193e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.141054242e-8
+ k1 = 5.952653582e-01 lk1 = -9.411969933e-9
+ k2 = -7.007272143e-02 lk2 = 8.434995606e-9
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 2.169351653e-01 ldsub = 4.203713551e-8
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.0054
+ cit = 0.0
+ voff = {-1.948584777e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -1.127067349e-8
+ nfactor = 1.941683786e+00 lnfactor = 2.237742136e-7
+ eta0 = -4.616715915e-01 leta0 = 4.531251049e-07 weta0 = 9.367506770e-23 peta0 = -9.887923813e-29
+ etab = -0.0003125
+ u0 = 2.386891122e-02 lu0 = 5.514072691e-11
+ ua = -1.285657146e-09 lua = 5.937146704e-17
+ ub = 1.885211294e-18 lub = -1.474075602e-25
+ uc = 7.885796353e-11 luc = -3.545029551e-17
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.618261931e+05 lvsat = 1.383556317e-2
+ a0 = 1.5
+ ags = 3.762869949e-01 lags = -1.698642534e-7
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = -5.168230143e-07 lb0 = 2.460780427e-13
+ b1 = 2.588712672e-08 lb1 = -1.232579297e-14
+ keta = 3.640521038e-02 lketa = -1.816720814e-08 pketa = -6.938893904e-30
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.429863183e+00 lpclm = -3.850497131e-7
+ pdiblc1 = 6.748458678e-01 lpdiblc1 = -8.340140914e-8
+ pdiblc2 = 1.013619654e-02 lpdiblc2 = -4.195314257e-09 wpdiblc2 = 6.938893904e-24
+ pdiblcb = -0.025
+ drout = 3.249506503e-01 ldrout = 3.214152972e-7
+ pscbe1 = 800000000.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = -5.127950400e-07 lalpha0 = 5.298417792e-13 walpha0 = 7.940933881e-29
+ alpha1 = 0.85
+ beta0 = 1.220304672e+01 lbeta0 = 1.617411747e-6
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -2.866014421e-01 lkt1 = -9.151194823e-9
+ kt2 = -4.153609621e-03 lkt2 = -2.177287003e-8
+ at = 2.537953600e+05 lat = -1.208411075e-1
+ ute = 9.716893932e-03 lute = -7.114517882e-7
+ ua1 = 3.923378182e-09 lua1 = -1.687764798e-15
+ ub1 = -2.711103396e-18 lub1 = 1.316087658e-24
+ uc1 = -8.391965094e-12 luc1 = 5.461861525e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -1.769019187e-03 ltvoff = -1.230720203e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.75e-6
+ sbref = 1.74e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.177 nmos
* Model Flag Parameters
+ lmin = 2.5e-07 lmax = 5.0e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {6.620950137e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = -4.816154384e-8
+ k1 = 2.755733038e-01 lk1 = 1.428049261e-7
+ k2 = 3.076911962e-02 lk2 = -3.957943522e-8
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 1.711988033e-02 ldsub = 1.371763860e-7
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 8.428413312e-03 lcdscd = -1.441936601e-9
+ cit = 0.0
+ voff = {-1.316296961e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = -4.137617264e-8
+ nfactor = 2.785225057e+00 lnfactor = -1.778661529e-7
+ eta0 = 9.332265600e-01 leta0 = -2.110361214e-7
+ etab = 3.920295691e-02 letab = -1.881473159e-08 wetab = 8.673617380e-25 petab = 1.192622390e-30
+ u0 = 2.353988335e-02 lu0 = 2.118027424e-10
+ ua = -1.157278411e-09 lua = -1.754270060e-18
+ ub = 1.248790162e-18 lub = 1.556154518e-25
+ uc = -7.434141045e-11 luc = 3.749344162e-17 wuc = -1.292469707e-32 puc = 9.693522803e-39
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 1.960511362e+05 lvsat = -2.460164352e-3
+ a0 = 1.5
+ ags = -1.093481875e+00 lags = 5.299456173e-07 wags = -8.326672685e-23 pags = 3.122502257e-29
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = 5.851559299e-02 lketa = -2.869475727e-08 pketa = -8.673617380e-31
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.019180347e+00 lpclm = -1.895088305e-7
+ pdiblc1 = 6.287709955e-01 lpdiblc1 = -6.146350373e-8
+ pdiblc2 = -5.080122993e-03 lpdiblc2 = 3.049723259e-09 wpdiblc2 = 1.734723476e-24 ppdiblc2 = -8.673617380e-31
+ pdiblcb = 4.582196898e-02 lpdiblcb = -3.372088902e-08 ppdiblcb = 6.938893904e-30
+ drout = 1.449262890e+00 ldrout = -2.139102352e-7
+ pscbe1 = 8.077610961e+08 lpscbe1 = -3.695337236e+0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.096051930e-06 lalpha0 = -2.361881816e-13
+ alpha1 = 0.85
+ beta0 = 1.668545280e+01 lbeta0 = -5.168231544e-7
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -3.825811247e-01 lkt1 = 3.654818732e-8
+ kt2 = -6.887994141e-02 lkt2 = 9.045666681e-9
+ at = -3.954710419e+04 lat = 1.882980000e-2
+ ute = -1.670350048e+00 lute = 8.848856547e-8
+ ua1 = 7.427581467e-10 lua1 = -1.733570974e-16
+ ub1 = -5.392589593e-19 lub1 = 2.819943349e-25 wub1 = 9.629649722e-41 pub1 = -3.611118646e-47
+ uc1 = 6.935515490e-11 luc1 = 1.760041252e-17
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.173720066e-03 ltvoff = 5.457566373e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.178 nmos
* Model Flag Parameters
+ lmin = 1.8e-07 lmax = 2.5e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {0.449119+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))}
+ k1 = 0.90707349
+ k2 = -0.1442558
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 0.62373
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-0.3146+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))}
+ nfactor = 1.99868
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 0.0244765
+ ua = -1.165036e-9
+ ub = 1.93694e-18
+ uc = 9.1459e-11
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 185172.0
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -0.068376
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 0.18115
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 5.16e-8
+ alpha1 = 0.85
+ beta0 = 14.4
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -0.22096074
+ kt2 = -0.028878939
+ at = 43720.487
+ ute = -1.2790432
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -0.00076032
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.1e-6
+ sbref = 1.1e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
* Well Proximity Effect Parameters
.model sky130_fd_pr__nfet_01v8.179 nmos
* Model Flag Parameters
+ lmin = 1.5e-07 lmax = 1.8e-07 wmin = 3.6e-07 wmax = 3.9e-7
+ level = 54.0
+ version = 4.5
+ binunit = 2.0
+ mobmod = 0.0
+ capmod = 2.0
+ igcmod = 0.0
+ igbmod = 0.0
+ geomod = 0.0
+ diomod = 1.0
+ rdsmod = 0.0
+ rbodymod = 1.0
+ rgatemod = 0.0
+ permod = 1.0
+ acnqsmod = 0.0
+ trnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ tempmod = 0.0
* Process Parameters
+ toxe = {4.148e-09+MC_MM_SWITCH*(4.148e-9*1.0*(sky130_fd_pr__nfet_01v8__toxe_slope/sqrt(1)))}
+ toxm = 4.148e-9
+ dtox = 0.0
+ epsrox = 3.9
+ xj = 1.5e-7
+ ngate = 1.0e+23
+ ndep = 1.7e+17
+ nsd = 1.0e+20
+ rsh = 1.0
+ rshg = 0.1
* Basic Model Parameters
+ wint = 2.1859e-8
+ lint = 1.1932e-8
+ vth0 = {-2.725906643e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__vth0_slope/sqrt(1))} lvth0 = 1.126848601e-07 wvth0 = 3.774853372e-07 pvth0 = -5.893905061e-14
+ k1 = 0.90707349
+ k2 = -4.780051754e-01 lk2 = 5.211029248e-08 wk2 = 1.485854542e-07 pk2 = -2.319953847e-14
+ k3 = 2.0
+ k3b = 0.54
+ w0 = 0.0
+ dvt0 = 0.0
+ dvt1 = 0.53
+ dvt2 = -0.032
+ dvt0w = -3.58
+ dvt1w = 1670600.0
+ dvt2w = 0.068
+ dsub = 3.327233912e+00 ldsub = -4.221142868e-07 wdsub = -1.017279859e-06 pdsub = 1.588340081e-13
+ minv = 0.0
+ voffl = 5.8197729e-9
+ lpe0 = 1.0325e-7
+ lpeb = -7.082e-8
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
+ phin = 0.0
+ cdsc = 0.0
+ cdscb = 0.0
+ cdscd = 0.002052
+ cit = 0.0
+ voff = {-7.647793840e-01+MC_MM_SWITCH*(sky130_fd_pr__nfet_01v8__voff_slope/sqrt(1))} lvoff = 7.028920830e-8
+ nfactor = -3.213434603e+00 lnfactor = 8.137987257e-07 wnfactor = 2.475245621e-07 pnfactor = -3.864749502e-14
+ eta0 = 0.0
+ etab = -0.043998
+ u0 = 8.608557677e-02 lu0 = -9.619394811e-09 wu0 = -4.705922369e-08 pu0 = 7.347638951e-15
+ ua = -1.393966070e-09 lua = 3.574422544e-17 wua = 1.398486904e-16 pua = -2.183541512e-23
+ ub = 6.496924862e-18 lub = -7.119777965e-25 wub = -2.980183442e-24 pub = 4.653139219e-31
+ uc = -1.261952913e-10 luc = 3.398367043e-17 wuc = 1.186133774e-16 puc = -1.851981829e-23
+ ud = 0.0
+ up = 0.0
+ lp = 1.0
+ eu = 1.67
+ vtl = 0.0
+ xn = 3.0
+ vsat = 3.539574068e+05 lvsat = -2.635347827e-02 wvsat = -8.318022480e-02 pvsat = 1.298742758e-8
+ a0 = 1.5
+ ags = 1.25
+ a1 = 0.0
+ a2 = 0.42385546
+ b0 = 0.0
+ b1 = 0.0
+ keta = -1.038255847e+00 lketa = 1.514331597e-07 wketa = 4.029564638e-07 pketa = -6.291601043e-14
+ dwg = 0.0
+ dwb = 0.0
+ pclm = 1.737607849e-02 lpclm = 2.557100501e-08 wpclm = 1.207637111e-07 ppclm = -1.885556280e-14
+ pdiblc1 = 0.35697215
+ pdiblc2 = 0.0084061121
+ pdiblcb = -0.10329577
+ drout = 0.50332666
+ pscbe1 = 791419880.0
+ pscbe2 = 1.0e-12
+ pvag = 0.0
+ delta = 0.01
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
+ lambda = 0.0
+ lc = 5.0e-9
* Parameters FOR Asymmetric AND Bias-Dependent RDS Model
+ rdsw = 65.968
+ rsw = 0.0
+ rdw = 0.0
+ rdswmin = 0.0
+ rdwmin = 0.0
+ rswmin = 0.0
+ prwb = 0.0
+ prwg = 0.021507
+ wr = 1.0
* Impact Ionization Current Model Parameters
+ alpha0 = 1.424179200e-07 lalpha0 = -1.417994676e-14 walpha0 = 2.191742220e-22 palpha0 = -3.422097810e-29
+ alpha1 = 0.85
+ beta0 = 1.671249334e+01 lbeta0 = -3.610634598e-07 wbeta0 = 3.836930773e-17 pbeta0 = -5.989875262e-24
* Gidl Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* Gate Dielectric Tunneling Current Model Parameters
+ toxref = 4.148e-9
+ dlcig = 0.0
+ aigbacc = 1.0
+ bigbacc = 0.0
+ cigbacc = 0.0
+ nigbacc = 0.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 0.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ nigc = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ vfbsdoff = 0.0
* Charge AND Capacitance Model Parameters
+ dlc = 9.87909e-9
+ dwc = 0.0
+ xpart = 0.0
+ cgso = 2.449068e-10
+ cgdo = 2.449068e-10
+ cgbo = 1.0e-13
+ cgdl = 0.0
+ cgsl = 0.0
+ clc = 1.0e-7
+ cle = 0.6
+ cf = 1.4067e-12
+ ckappas = 0.6
+ vfbcv = -1.0
+ acde = 0.4
+ moin = 6.9
+ noff = 3.4037
+ voffcv = -0.17287
* High-Speed/RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* Flicker AND Thermal Noise Model Parameters
+ ef = 0.84
+ noia = 2.5e+42
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ ntnoi = 1.0
+ lintnoi = -1.0e-7
+ af = 1.0
+ kf = 0.0
+ tnoia = 15000000.0
+ tnoib = 9900000.0
+ rnoia = 0.94
+ rnoib = 0.26
* Layout-Dependent Parasitics Model Parameters
+ xl = 0.0
+ xw = 0.0
+ dmcg = 0.0
+ dmdg = 0.0
+ dmcgt = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Asymmetric Source/Drain Junction Diode Model Parameters
+ jss = 0.00275
+ jsws = 6.0e-10
+ ijthsfwd = 0.1
+ ijthsrev = 0.1
+ bvs = 11.7
+ xjbvs = 1.0
+ pbs = 0.729
+ cjs = 0.001339749237
+ mjs = 0.44
+ pbsws = 0.2
+ cjsws = 3.67354204e-11
+ mjsws = 0.0009
+ pbswgs = 0.95578
+ cjswgs = 2.38232788e-10
+ mjswgs = 0.8
* Temperature Dependence Parameters
+ tnom = 30.0
+ kt1 = -1.368700733e-01 lkt1 = -1.312958033e-08 wkt1 = -8.156852971e-17 pkt1 = 1.273581240e-23
+ kt2 = -0.028878939
+ at = 1.675153666e+03 lat = 6.564790165e-03 wat = -2.587959170e-11 pat = 4.040746717e-18
+ ute = -9.418347116e-01 lute = -5.265038454e-08 wute = -2.218108973e-07 pute = 3.463266627e-14
+ ua1 = -2.3847336e-11
+ ub1 = 7.0775317e-19
+ uc1 = 1.4718625e-10
+ kt1l = 0.0
+ prt = 0.0
+ tvoff = -3.957110784e-03 ltvoff = 4.991341259e-10
+ njs = 1.2928
+ tpb = 0.0012287
+ tcj = 0.000792
+ tpbsw = 0.0
+ tcjsw = 1.0e-5
+ tpbswg = 0.0
+ tcjswg = 0.0
+ xtis = 2.0
+ tvfbsdoff = 0.0
* DW AND DL Parameters
+ ll = 0.0
+ wl = 0.0
+ lln = 1.0
+ wln = 1.0
+ lw = 0.0
+ ww = 0.0
+ lwn = 1.0
+ wwn = 1.0
+ lwl = 0.0
+ wwl = 0.0
+ llc = 0.0
+ wlc = 0.0
+ lwc = 0.0
+ wwc = 0.0
+ lwlc = 0.0
+ wwlc = 0.0
* Stress Parameters
+ saref = 1.04e-6
+ sbref = 1.04e-6
+ kvth0 = 9.8e-9
+ lkvth0 = 0.0
+ wkvth0 = 2.0e-7
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ wlod = 0.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = -2.7e-8
+ lku0 = 0.0
+ wku0 = 0.0
+ pku0 = 0.0
+ tku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = 0.2
+ steta0 = 0.0
.ends sky130_fd_pr__nfet_01v8
* Well Proximity Effect Parameters
