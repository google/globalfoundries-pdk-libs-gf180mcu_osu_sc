

.option scale=0.05u

.subckt gf180mcu_osu_sc_9T_xnor2_1 A Y B
X0 a_42_70 a_9_19 VDD VDD pmos_3p3 w=34 l=6
X1 Y a_49_14 a_42_70 VDD pmos_3p3 w=34 l=6
X2 a_49_14 B VDD VDD pmos_3p3 w=34 l=6
X3 GND A a_9_19 GND nmos_3p3 w=17 l=6
X4 VDD A a_9_19 VDD pmos_3p3 w=34 l=6
X5 a_78_19 a_9_19 Y GND nmos_3p3 w=17 l=6
X6 GND B a_78_19 GND nmos_3p3 w=17 l=6
X7 a_78_70 A Y VDD pmos_3p3 w=34 l=6
X8 a_42_19 A GND GND nmos_3p3 w=17 l=6
X9 VDD B a_78_70 VDD pmos_3p3 w=34 l=6
X10 Y a_49_14 a_42_19 GND nmos_3p3 w=17 l=6
X11 a_49_14 B GND GND nmos_3p3 w=17 l=6
.ends

