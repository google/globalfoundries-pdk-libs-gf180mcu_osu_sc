# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__clkbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__clkbuf_1 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 1.4 3.5 1.75 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 1.4 0 1.75 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.85 1.55 3.15 ;
      LAYER MET2 ;
        RECT 1.05 2.85 1.55 3.15 ;
        RECT 1.1 2.8 1.5 3.2 ;
      LAYER VIA12 ;
        RECT 1.17 2.87 1.43 3.13 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 1.5 2.75 1.8 ;
        RECT 2.35 0.95 2.6 1.8 ;
        RECT 2.25 3.5 2.75 3.8 ;
        RECT 2.35 3.5 2.6 5.2 ;
      LAYER MET2 ;
        RECT 2.25 3.45 2.75 3.85 ;
        RECT 2.25 1.45 2.75 1.85 ;
        RECT 2.35 1.45 2.65 3.85 ;
      LAYER VIA12 ;
        RECT 2.37 3.52 2.63 3.78 ;
        RECT 2.37 1.52 2.63 1.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.15 2.2 2.45 ;
  END
END gf180mcu_osu_sc_gp9t3v3__clkbuf_1
