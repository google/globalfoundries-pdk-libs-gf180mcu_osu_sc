# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__dff_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__dff_1 0 0 ;
  SIZE 14.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 14.5 6.15 ;
        RECT 12.85 4.05 13.1 6.15 ;
        RECT 10.4 3.5 10.65 6.15 ;
        RECT 8.6 4.75 8.85 6.15 ;
        RECT 5 4.1 5.25 6.15 ;
        RECT 1.4 4.75 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 14.5 0.6 ;
        RECT 12.85 0 13.1 1.6 ;
        RECT 10.4 0 10.65 1.4 ;
        RECT 8.6 0 8.85 1.5 ;
        RECT 5 0 5.25 1.4 ;
        RECT 1.4 0 1.65 1.5 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 2.5 3 9.4 3.25 ;
        RECT 2.5 3 8.95 3.3 ;
        RECT 5.95 1.95 6.45 2.25 ;
        RECT 6.05 1.95 6.35 3.3 ;
        RECT 3.8 2 4.3 2.3 ;
        RECT 3.9 2 4.2 3.3 ;
      LAYER MET2 ;
        RECT 9 2.85 9.5 3.15 ;
        RECT 9.05 2.8 9.45 3.2 ;
      LAYER VIA12 ;
        RECT 9.12 2.87 9.38 3.13 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 2.85 2.25 3.15 ;
      LAYER MET2 ;
        RECT 1.7 2.85 2.3 3.15 ;
        RECT 1.75 2.8 2.25 3.2 ;
      LAYER VIA12 ;
        RECT 1.87 2.87 2.13 3.13 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 13.7 4.15 14.25 4.5 ;
        RECT 13.7 4.1 14.2 4.5 ;
        RECT 13.7 0.95 13.95 5.2 ;
      LAYER MET2 ;
        RECT 13.75 4.15 14.25 4.45 ;
        RECT 13.8 4.1 14.2 4.5 ;
      LAYER VIA12 ;
        RECT 13.87 4.17 14.13 4.43 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12 3.5 13.45 3.8 ;
        RECT 13.05 1.85 13.35 3.8 ;
        RECT 12 1.85 13.35 2.1 ;
        RECT 12 3.5 12.25 5.2 ;
        RECT 12 0.95 12.25 2.1 ;
      LAYER MET2 ;
        RECT 12.95 3.5 13.45 3.8 ;
        RECT 13 3.45 13.4 3.85 ;
      LAYER VIA12 ;
        RECT 13.07 3.52 13.33 3.78 ;
    END
  END QN
  OBS
    LAYER MET2 ;
      RECT 8.1 4.15 8.5 4.55 ;
      RECT 8.05 4.2 11.45 4.5 ;
      RECT 11.15 2.55 11.45 4.5 ;
      RECT 8.15 2.15 8.45 4.55 ;
      RECT 12.2 2.5 12.6 2.9 ;
      RECT 11.15 2.55 12.65 2.85 ;
      RECT 8.1 2.15 8.5 2.55 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 6.4 0.9 6.7 4.6 ;
      RECT 6.35 4.15 6.75 4.55 ;
      RECT 10.55 1.6 10.95 2 ;
      RECT 10.2 1.65 11 1.95 ;
      RECT 6.35 1.3 6.75 1.7 ;
      RECT 6.4 0.9 6.75 1.7 ;
      RECT 6.3 1.35 6.75 1.65 ;
      RECT 10.2 1.6 10.95 1.95 ;
      RECT 10.2 0.9 10.5 1.95 ;
      RECT 6.4 0.9 10.5 1.2 ;
      RECT 2.8 4.9 7.55 5.2 ;
      RECT 7.25 1.5 7.55 5.2 ;
      RECT 2.8 1.95 3.1 5.2 ;
      RECT 2.75 1.95 3.2 2.35 ;
      RECT 2.7 2 3.2 2.3 ;
      RECT 9.4 1.5 9.8 1.9 ;
      RECT 7.2 1.5 7.6 1.9 ;
      RECT 7.15 1.55 9.9 1.85 ;
      RECT 4.65 1.95 5.05 2.35 ;
      RECT 0.45 1.95 0.85 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 0.4 2 0.9 2.3 ;
      RECT 4.7 1.05 5 2.35 ;
      RECT 0.5 1.05 0.8 2.35 ;
      RECT 0.5 1.05 5 1.35 ;
    LAYER VIA12 ;
      RECT 12.27 2.57 12.53 2.83 ;
      RECT 10.62 1.67 10.88 1.93 ;
      RECT 9.47 1.57 9.73 1.83 ;
      RECT 8.17 2.22 8.43 2.48 ;
      RECT 8.17 4.22 8.43 4.48 ;
      RECT 7.27 1.57 7.53 1.83 ;
      RECT 6.42 1.37 6.68 1.63 ;
      RECT 6.42 4.22 6.68 4.48 ;
      RECT 4.72 2.02 4.98 2.28 ;
      RECT 2.82 2.02 3.08 2.28 ;
      RECT 0.52 2.02 0.78 2.28 ;
    LAYER MET1 ;
      RECT 11.25 0.95 11.5 5.2 ;
      RECT 11.25 2.55 12.65 2.85 ;
      RECT 10.6 1.65 10.9 2.95 ;
      RECT 10.5 1.65 11 1.95 ;
      RECT 9.45 3.5 9.7 5.2 ;
      RECT 9.45 3.5 10 3.75 ;
      RECT 9.75 2.2 10 3.75 ;
      RECT 9.45 1.45 9.75 2.5 ;
      RECT 9.45 0.95 9.7 2.5 ;
      RECT 8.05 4.2 8.55 4.5 ;
      RECT 8.15 4.1 8.45 4.5 ;
      RECT 6.95 1.9 7.25 2.4 ;
      RECT 6.9 2 7.55 2.3 ;
      RECT 7.25 1.45 7.55 2.3 ;
      RECT 6.3 1.4 6.95 1.65 ;
      RECT 6.4 0.95 6.95 1.65 ;
      RECT 6.4 4.2 6.95 5.2 ;
      RECT 6.4 4.1 6.7 5.2 ;
      RECT 4.7 2 5 2.35 ;
      RECT 4.6 2 5.1 2.3 ;
      RECT 3.3 4.2 3.85 5.2 ;
      RECT 1.05 4.2 3.85 4.5 ;
      RECT 1.05 1.8 1.35 4.5 ;
      RECT 1.05 3 1.45 3.3 ;
      RECT 1.05 1.8 2.25 2.05 ;
      RECT 2 1.4 2.25 2.05 ;
      RECT 2 1.4 3.85 1.65 ;
      RECT 3.3 0.95 3.85 1.65 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.5 1.9 0.8 2.35 ;
      RECT 0.4 2 0.8 2.3 ;
      RECT 8.05 2.2 8.55 2.5 ;
      RECT 2.7 2 3.2 2.3 ;
  END
END gf180mcu_osu_sc_gp9t3v3__dff_1
