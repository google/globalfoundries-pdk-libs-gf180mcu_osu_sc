magic
tech gf180mcuC
timestamp 1660079376
<< error_p >>
rect 16 97 18 159
<< nwell >>
rect 0 97 16 159
<< metal1 >>
rect 0 147 16 159
rect 0 -3 16 9
<< labels >>
rlabel metal1 7 154 7 154 5 VDD
rlabel metal1 6 2 6 2 1 GND
<< end >>
