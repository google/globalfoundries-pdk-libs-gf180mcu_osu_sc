# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__oai22_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai22_1 0 0 ;
  SIZE 5.5 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 5.5 6.35 ;
        RECT 3.6 3.6 3.85 6.35 ;
        RECT 0.65 3.6 0.9 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.5 0.7 ;
        RECT 1.35 0 1.6 1.55 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 2.3 1.2 2.6 ;
      LAYER Metal2 ;
        RECT 0.7 2.25 1.2 2.65 ;
      LAYER Via1 ;
        RECT 0.82 2.32 1.08 2.58 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.65 2.3 2.15 2.6 ;
      LAYER Metal2 ;
        RECT 1.65 2.25 2.15 2.65 ;
      LAYER Via1 ;
        RECT 1.77 2.32 2.03 2.58 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.55 2.3 3.05 2.6 ;
      LAYER Metal2 ;
        RECT 2.55 2.25 3.05 2.65 ;
      LAYER Via1 ;
        RECT 2.67 2.32 2.93 2.58 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.35 2.3 3.85 2.6 ;
      LAYER Metal2 ;
        RECT 3.35 2.25 3.85 2.65 ;
      LAYER Via1 ;
        RECT 3.47 2.32 3.73 2.58 ;
    END
  END B1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4.5 0.95 5 1.25 ;
        RECT 2.1 2.85 4.9 3.15 ;
        RECT 4.6 0.95 4.9 3.15 ;
        RECT 2.1 2.85 2.45 5.3 ;
        RECT 3.05 0.95 3.55 1.3 ;
        RECT 3.15 0.95 3.4 1.55 ;
      LAYER Metal2 ;
        RECT 3.05 0.95 5 1.25 ;
        RECT 4.55 0.9 4.95 1.3 ;
        RECT 3.05 0.9 3.55 1.3 ;
      LAYER Via1 ;
        RECT 3.17 0.97 3.43 1.23 ;
        RECT 4.62 0.97 4.88 1.23 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 0.5 1.8 4.25 2.05 ;
      RECT 4 1.05 4.25 2.05 ;
      RECT 2.2 1.05 2.55 2.05 ;
      RECT 0.5 1.05 0.75 2.05 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai22_1
