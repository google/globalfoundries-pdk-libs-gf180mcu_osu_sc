# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifup 0 0 ;
  SIZE 7.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 2.3 8.1 ;
        RECT 0.55 5.45 0.85 8.1 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.9 7.5 7.8 8.1 ;
        RECT 6.05 5.45 6.35 8.1 ;
        RECT 4.35 5.45 4.65 8.1 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 7.8 0.6 ;
        RECT 6.05 0 6.35 1.8 ;
        RECT 4.35 0 4.65 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4 2.2 4.5 2.5 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 4 2.15 4.5 2.55 ;
        RECT 0.6 2.2 4.5 2.5 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
        RECT 4.12 2.22 4.38 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 6.9 4.15 7.3 4.45 ;
        RECT 6.95 0.95 7.25 7.15 ;
      LAYER MET2 ;
        RECT 6.85 4.1 7.35 4.5 ;
      LAYER VIA12 ;
        RECT 6.97 4.17 7.23 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 6.1 4.75 6.6 5.15 ;
      RECT 4.55 4.75 4.95 5.15 ;
      RECT 4.5 4.8 6.6 5.1 ;
      RECT 4.5 2.85 5 3.25 ;
      RECT 1.35 2.85 1.85 3.25 ;
      RECT 1.35 2.9 5 3.2 ;
    LAYER VIA12 ;
      RECT 6.22 4.82 6.48 5.08 ;
      RECT 4.62 2.92 4.88 3.18 ;
      RECT 4.62 4.82 4.88 5.08 ;
      RECT 1.47 2.92 1.73 3.18 ;
    LAYER MET1 ;
      RECT 5.25 0.95 5.55 7.15 ;
      RECT 4.8 4 5.55 4.45 ;
      RECT 3.45 0.95 3.75 7.15 ;
      RECT 4.55 4.75 5 5.2 ;
      RECT 3.45 4.8 5 5.1 ;
      RECT 1.45 0.95 1.75 7.15 ;
      RECT 1.35 2.9 1.85 3.2 ;
      RECT 6.1 4.8 6.6 5.1 ;
      RECT 4.5 2.9 5 3.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifup
