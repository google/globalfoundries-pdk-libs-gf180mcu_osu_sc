magic
tech gf180mcuC
timestamp 1661529368
<< nwell >>
rect 0 97 290 159
<< nmos >>
rect 19 55 25 72
rect 36 55 42 72
rect 57 55 63 72
rect 80 55 86 72
rect 91 55 97 72
rect 108 55 114 72
rect 119 55 125 72
rect 142 55 148 72
rect 163 55 169 72
rect 180 55 186 72
rect 216 55 222 72
rect 248 55 254 72
rect 265 55 271 72
<< pmos >>
rect 19 106 25 140
rect 36 106 42 140
rect 57 106 63 140
rect 80 106 86 140
rect 91 106 97 140
rect 108 106 114 140
rect 119 106 125 140
rect 142 106 148 140
rect 163 106 169 140
rect 180 106 186 140
rect 216 106 222 140
rect 248 106 254 140
rect 265 106 271 140
<< ndiff >>
rect 9 70 19 72
rect 9 57 11 70
rect 16 57 19 70
rect 9 55 19 57
rect 25 63 36 72
rect 25 57 28 63
rect 33 57 36 63
rect 25 55 36 57
rect 42 55 57 72
rect 63 63 80 72
rect 63 57 66 63
rect 77 57 80 63
rect 63 55 80 57
rect 86 55 91 72
rect 97 62 108 72
rect 97 57 100 62
rect 105 57 108 62
rect 97 55 108 57
rect 114 55 119 72
rect 125 62 142 72
rect 125 57 128 62
rect 139 57 142 62
rect 125 55 142 57
rect 148 55 163 72
rect 169 63 180 72
rect 169 57 172 63
rect 177 57 180 63
rect 169 55 180 57
rect 186 62 196 72
rect 186 57 189 62
rect 194 57 196 62
rect 186 55 196 57
rect 206 62 216 72
rect 206 57 208 62
rect 213 57 216 62
rect 206 55 216 57
rect 222 70 232 72
rect 222 57 225 70
rect 230 57 232 70
rect 222 55 232 57
rect 238 70 248 72
rect 238 57 240 70
rect 245 57 248 70
rect 238 55 248 57
rect 254 66 265 72
rect 254 57 257 66
rect 262 57 265 66
rect 254 55 265 57
rect 271 70 281 72
rect 271 57 274 70
rect 279 57 281 70
rect 271 55 281 57
<< pdiff >>
rect 9 138 19 140
rect 9 108 11 138
rect 16 108 19 138
rect 9 106 19 108
rect 25 138 36 140
rect 25 133 28 138
rect 33 133 36 138
rect 25 106 36 133
rect 42 106 57 140
rect 63 138 80 140
rect 63 122 66 138
rect 77 122 80 138
rect 63 106 80 122
rect 86 106 91 140
rect 97 138 108 140
rect 97 120 100 138
rect 105 120 108 138
rect 97 106 108 120
rect 114 106 119 140
rect 125 138 142 140
rect 125 122 128 138
rect 139 122 142 138
rect 125 106 142 122
rect 148 106 163 140
rect 169 138 180 140
rect 169 133 172 138
rect 177 133 180 138
rect 169 106 180 133
rect 186 138 196 140
rect 186 108 189 138
rect 194 108 196 138
rect 186 106 196 108
rect 206 138 216 140
rect 206 108 208 138
rect 213 108 216 138
rect 206 106 216 108
rect 222 138 232 140
rect 222 108 225 138
rect 230 108 232 138
rect 222 106 232 108
rect 238 138 248 140
rect 238 108 240 138
rect 245 108 248 138
rect 238 106 248 108
rect 254 138 265 140
rect 254 119 257 138
rect 262 119 265 138
rect 254 106 265 119
rect 271 138 281 140
rect 271 125 274 138
rect 279 125 281 138
rect 271 106 281 125
<< ndiffc >>
rect 11 57 16 70
rect 28 57 33 63
rect 66 57 77 63
rect 100 57 105 62
rect 128 57 139 62
rect 172 57 177 63
rect 189 57 194 62
rect 208 57 213 62
rect 225 57 230 70
rect 240 57 245 70
rect 257 57 262 66
rect 274 57 279 70
<< pdiffc >>
rect 11 108 16 138
rect 28 133 33 138
rect 66 122 77 138
rect 100 120 105 138
rect 128 122 139 138
rect 172 133 177 138
rect 189 108 194 138
rect 208 108 213 138
rect 225 108 230 138
rect 240 108 245 138
rect 257 119 262 138
rect 274 125 279 138
<< psubdiff >>
rect 9 46 18 48
rect 9 41 11 46
rect 16 41 18 46
rect 9 39 18 41
rect 33 46 42 48
rect 33 41 35 46
rect 40 41 42 46
rect 33 39 42 41
rect 57 46 66 48
rect 57 41 59 46
rect 64 41 66 46
rect 57 39 66 41
rect 81 46 90 48
rect 81 41 83 46
rect 88 41 90 46
rect 81 39 90 41
rect 105 46 114 48
rect 105 41 107 46
rect 112 41 114 46
rect 105 39 114 41
rect 129 46 138 48
rect 129 41 131 46
rect 136 41 138 46
rect 129 39 138 41
rect 153 46 162 48
rect 153 41 155 46
rect 160 41 162 46
rect 153 39 162 41
rect 177 46 186 48
rect 177 41 179 46
rect 184 41 186 46
rect 177 39 186 41
rect 201 46 210 48
rect 201 41 203 46
rect 208 41 210 46
rect 201 39 210 41
rect 225 46 234 48
rect 225 41 227 46
rect 232 41 234 46
rect 225 39 234 41
rect 249 46 258 48
rect 249 41 251 46
rect 256 41 258 46
rect 249 39 258 41
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
rect 81 154 90 156
rect 81 149 83 154
rect 88 149 90 154
rect 81 147 90 149
rect 105 154 114 156
rect 105 149 107 154
rect 112 149 114 154
rect 105 147 114 149
rect 129 154 138 156
rect 129 149 131 154
rect 136 149 138 154
rect 129 147 138 149
rect 153 154 162 156
rect 153 149 155 154
rect 160 149 162 154
rect 153 147 162 149
rect 177 154 186 156
rect 177 149 179 154
rect 184 149 186 154
rect 177 147 186 149
rect 201 154 210 156
rect 201 149 203 154
rect 208 149 210 154
rect 201 147 210 149
rect 225 154 234 156
rect 225 149 227 154
rect 232 149 234 154
rect 225 147 234 149
rect 249 154 258 156
rect 249 149 251 154
rect 256 149 258 154
rect 249 147 258 149
<< psubdiffcont >>
rect 11 41 16 46
rect 35 41 40 46
rect 59 41 64 46
rect 83 41 88 46
rect 107 41 112 46
rect 131 41 136 46
rect 155 41 160 46
rect 179 41 184 46
rect 203 41 208 46
rect 227 41 232 46
rect 251 41 256 46
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
rect 83 149 88 154
rect 107 149 112 154
rect 131 149 136 154
rect 155 149 160 154
rect 179 149 184 154
rect 203 149 208 154
rect 227 149 232 154
rect 251 149 256 154
<< polysilicon >>
rect 19 140 25 145
rect 36 140 42 145
rect 57 140 63 145
rect 80 140 86 145
rect 91 140 97 145
rect 108 140 114 145
rect 119 140 125 145
rect 142 140 148 145
rect 163 140 169 145
rect 180 140 186 145
rect 216 140 222 145
rect 248 140 254 145
rect 265 140 271 145
rect 19 104 25 106
rect 19 102 29 104
rect 19 96 21 102
rect 27 96 29 102
rect 36 101 42 106
rect 57 104 63 106
rect 50 102 63 104
rect 19 94 29 96
rect 34 99 45 101
rect 19 72 25 94
rect 34 93 37 99
rect 43 93 45 99
rect 50 97 53 102
rect 58 101 63 102
rect 58 97 60 101
rect 50 95 60 97
rect 80 93 86 106
rect 91 104 97 106
rect 108 104 114 106
rect 91 97 114 104
rect 34 91 45 93
rect 36 72 42 91
rect 65 88 86 93
rect 65 84 71 88
rect 53 82 71 84
rect 99 83 105 97
rect 119 93 125 106
rect 142 104 148 106
rect 142 102 154 104
rect 142 101 146 102
rect 144 96 146 101
rect 152 96 154 102
rect 144 94 154 96
rect 119 88 139 93
rect 163 88 169 106
rect 180 101 186 106
rect 180 99 190 101
rect 180 93 182 99
rect 188 93 190 99
rect 216 95 222 106
rect 248 95 254 106
rect 180 91 190 93
rect 210 93 222 95
rect 134 86 139 88
rect 161 86 171 88
rect 53 76 56 82
rect 62 76 71 82
rect 76 81 86 83
rect 76 76 78 81
rect 84 76 86 81
rect 53 74 65 76
rect 76 74 86 76
rect 57 72 63 74
rect 80 72 86 74
rect 91 82 105 83
rect 91 81 114 82
rect 91 76 94 81
rect 100 76 114 81
rect 91 74 114 76
rect 91 72 97 74
rect 108 72 114 74
rect 119 81 129 83
rect 119 76 121 81
rect 127 76 129 81
rect 134 82 148 86
rect 134 76 139 82
rect 145 76 148 82
rect 161 80 163 86
rect 169 80 171 86
rect 161 78 171 80
rect 119 74 129 76
rect 137 74 148 76
rect 119 72 125 74
rect 142 72 148 74
rect 163 72 169 78
rect 180 72 186 91
rect 210 87 212 93
rect 218 87 222 93
rect 210 85 222 87
rect 243 93 254 95
rect 243 87 245 93
rect 251 87 254 93
rect 265 88 271 106
rect 243 85 254 87
rect 216 72 222 85
rect 248 72 254 85
rect 259 86 271 88
rect 259 80 261 86
rect 267 80 271 86
rect 259 78 271 80
rect 265 72 271 78
rect 19 50 25 55
rect 36 50 42 55
rect 57 50 63 55
rect 80 50 86 55
rect 91 50 97 55
rect 108 50 114 55
rect 119 50 125 55
rect 142 50 148 55
rect 163 50 169 55
rect 180 50 186 55
rect 216 50 222 55
rect 248 50 254 55
rect 265 50 271 55
<< polycontact >>
rect 21 96 27 102
rect 37 93 43 99
rect 53 97 58 102
rect 146 96 152 102
rect 182 93 188 99
rect 56 76 62 82
rect 78 76 84 81
rect 94 76 100 81
rect 121 76 127 81
rect 139 76 145 82
rect 163 80 169 86
rect 212 87 218 93
rect 245 87 251 93
rect 261 80 267 86
<< metal1 >>
rect 0 154 290 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 83 154
rect 89 148 107 154
rect 113 148 131 154
rect 137 148 155 154
rect 161 148 179 154
rect 185 148 203 154
rect 209 148 227 154
rect 233 148 251 154
rect 257 148 290 154
rect 0 147 290 148
rect 11 138 16 140
rect 28 138 33 147
rect 28 131 33 133
rect 66 138 77 140
rect 11 83 16 108
rect 10 82 16 83
rect 8 76 10 82
rect 10 74 16 76
rect 11 70 16 74
rect 21 122 66 126
rect 21 120 77 122
rect 100 138 105 147
rect 21 102 27 120
rect 100 118 105 120
rect 128 138 139 140
rect 172 138 177 147
rect 172 131 177 133
rect 189 138 194 140
rect 134 120 139 122
rect 161 120 163 126
rect 169 120 171 126
rect 128 118 134 120
rect 163 118 169 120
rect 208 138 213 147
rect 194 108 200 111
rect 189 106 200 108
rect 208 106 213 108
rect 225 138 230 140
rect 27 96 29 102
rect 21 77 27 96
rect 35 93 37 99
rect 43 93 45 99
rect 50 97 53 102
rect 58 97 146 102
rect 50 96 146 97
rect 152 101 179 102
rect 152 99 188 101
rect 152 96 182 99
rect 78 82 84 96
rect 94 82 100 83
rect 21 72 45 77
rect 54 76 56 82
rect 62 76 64 82
rect 76 81 86 82
rect 76 76 78 81
rect 84 76 86 81
rect 92 76 94 82
rect 100 76 102 82
rect 121 81 127 96
rect 180 93 182 96
rect 188 93 190 99
rect 195 86 200 106
rect 139 82 145 84
rect 119 76 121 81
rect 127 76 129 81
rect 138 76 139 82
rect 145 76 151 82
rect 161 80 163 86
rect 169 80 171 86
rect 189 80 200 86
rect 212 93 218 95
rect 119 75 129 76
rect 139 74 151 76
rect 40 69 45 72
rect 145 73 151 74
rect 11 55 16 57
rect 28 63 33 66
rect 40 64 77 69
rect 126 64 128 69
rect 28 48 33 57
rect 66 63 77 64
rect 66 55 77 57
rect 100 62 105 64
rect 100 48 105 57
rect 134 63 139 69
rect 145 65 151 67
rect 189 73 195 80
rect 212 75 218 87
rect 225 93 230 108
rect 240 138 245 140
rect 257 138 262 147
rect 257 117 262 119
rect 274 138 279 140
rect 279 125 285 126
rect 274 119 277 125
rect 283 119 285 125
rect 274 118 284 119
rect 245 108 261 112
rect 240 106 261 108
rect 267 106 269 112
rect 225 87 245 93
rect 251 87 253 93
rect 210 69 212 75
rect 218 69 220 75
rect 225 70 230 87
rect 261 86 267 106
rect 261 78 267 80
rect 128 62 139 63
rect 128 55 139 57
rect 172 63 177 66
rect 172 48 177 57
rect 189 65 195 67
rect 189 62 194 65
rect 189 55 194 57
rect 208 62 213 64
rect 208 48 213 57
rect 225 55 230 57
rect 240 73 267 78
rect 240 70 245 73
rect 274 70 279 118
rect 240 55 245 57
rect 257 66 262 68
rect 257 48 262 57
rect 274 55 279 57
rect 0 47 290 48
rect 0 41 11 47
rect 17 41 35 47
rect 41 41 59 47
rect 65 41 83 47
rect 89 41 107 47
rect 113 41 131 47
rect 137 41 155 47
rect 161 41 179 47
rect 185 41 203 47
rect 209 41 227 47
rect 233 41 251 47
rect 257 41 290 47
rect 0 36 290 41
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 83 149 88 154
rect 88 149 89 154
rect 83 148 89 149
rect 107 149 112 154
rect 112 149 113 154
rect 107 148 113 149
rect 131 149 136 154
rect 136 149 137 154
rect 131 148 137 149
rect 155 149 160 154
rect 160 149 161 154
rect 155 148 161 149
rect 179 149 184 154
rect 184 149 185 154
rect 179 148 185 149
rect 203 149 208 154
rect 208 149 209 154
rect 203 148 209 149
rect 227 149 232 154
rect 232 149 233 154
rect 227 148 233 149
rect 251 149 256 154
rect 256 149 257 154
rect 251 148 257 149
rect 10 76 16 82
rect 128 122 134 126
rect 128 120 134 122
rect 163 120 169 126
rect 37 93 43 99
rect 56 76 62 82
rect 94 81 100 82
rect 94 76 100 81
rect 182 93 188 99
rect 163 80 169 86
rect 128 63 134 69
rect 145 67 151 73
rect 277 119 283 125
rect 261 106 267 112
rect 245 87 251 93
rect 189 67 195 73
rect 212 69 218 75
rect 11 46 17 47
rect 11 41 16 46
rect 16 41 17 46
rect 35 46 41 47
rect 35 41 40 46
rect 40 41 41 46
rect 59 46 65 47
rect 59 41 64 46
rect 64 41 65 46
rect 83 46 89 47
rect 83 41 88 46
rect 88 41 89 46
rect 107 46 113 47
rect 107 41 112 46
rect 112 41 113 46
rect 131 46 137 47
rect 131 41 136 46
rect 136 41 137 46
rect 155 46 161 47
rect 155 41 160 46
rect 160 41 161 46
rect 179 46 185 47
rect 179 41 184 46
rect 184 41 185 46
rect 203 46 209 47
rect 203 41 208 46
rect 208 41 209 46
rect 227 46 233 47
rect 227 41 232 46
rect 232 41 233 46
rect 251 46 257 47
rect 251 41 256 46
rect 256 41 257 46
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 130 154 138 155
rect 154 154 162 155
rect 178 154 186 155
rect 202 154 210 155
rect 226 154 234 155
rect 250 154 258 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 81 148 83 154
rect 89 148 91 154
rect 105 148 107 154
rect 113 148 115 154
rect 129 148 131 154
rect 137 148 139 154
rect 153 148 155 154
rect 161 148 163 154
rect 177 148 179 154
rect 185 148 187 154
rect 201 148 203 154
rect 209 148 211 154
rect 225 148 227 154
rect 233 148 235 154
rect 249 148 251 154
rect 257 148 259 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 130 147 138 148
rect 154 147 162 148
rect 178 147 186 148
rect 202 147 210 148
rect 226 147 234 148
rect 250 147 258 148
rect 56 134 151 140
rect 35 99 45 100
rect 34 93 37 99
rect 43 93 46 99
rect 35 92 45 93
rect 56 83 62 134
rect 128 127 134 128
rect 127 126 135 127
rect 127 120 128 126
rect 134 120 135 126
rect 127 119 135 120
rect 9 82 17 83
rect 55 82 64 83
rect 93 82 101 83
rect 8 76 10 82
rect 16 76 18 82
rect 54 76 56 82
rect 62 76 64 82
rect 92 76 94 82
rect 100 76 102 82
rect 9 75 17 76
rect 55 75 64 76
rect 93 75 101 76
rect 10 63 16 75
rect 94 63 100 75
rect 128 70 134 119
rect 145 74 151 134
rect 162 126 170 127
rect 161 120 163 126
rect 169 120 229 126
rect 276 125 284 126
rect 162 119 170 120
rect 163 87 169 119
rect 181 99 189 100
rect 180 93 182 99
rect 188 93 190 99
rect 223 93 229 120
rect 275 119 277 125
rect 283 119 285 125
rect 276 118 284 119
rect 260 112 268 113
rect 259 106 261 112
rect 267 106 269 112
rect 260 105 268 106
rect 244 93 252 94
rect 181 92 189 93
rect 223 87 245 93
rect 251 87 253 93
rect 162 86 170 87
rect 244 86 252 87
rect 161 80 163 86
rect 169 80 171 86
rect 162 79 170 80
rect 211 75 219 76
rect 144 73 152 74
rect 188 73 196 74
rect 127 69 135 70
rect 126 63 128 69
rect 134 63 135 69
rect 143 67 145 73
rect 151 67 189 73
rect 195 67 198 73
rect 204 69 212 75
rect 218 69 220 75
rect 204 68 219 69
rect 144 66 152 67
rect 188 66 196 67
rect 10 57 100 63
rect 127 62 135 63
rect 128 60 135 62
rect 204 60 210 68
rect 128 54 210 60
rect 10 47 18 48
rect 34 47 42 48
rect 58 47 66 48
rect 82 47 90 48
rect 106 47 114 48
rect 130 47 138 48
rect 154 47 162 48
rect 178 47 186 48
rect 202 47 210 48
rect 226 47 234 48
rect 250 47 258 48
rect 9 41 11 47
rect 17 41 19 47
rect 33 41 35 47
rect 41 41 43 47
rect 57 41 59 47
rect 65 41 67 47
rect 81 41 83 47
rect 89 41 91 47
rect 105 41 107 47
rect 113 41 115 47
rect 129 41 131 47
rect 137 41 139 47
rect 153 41 155 47
rect 161 41 163 47
rect 177 41 179 47
rect 185 41 187 47
rect 201 41 203 47
rect 209 41 211 47
rect 225 41 227 47
rect 233 41 235 47
rect 249 41 251 47
rect 257 41 259 47
rect 10 40 18 41
rect 34 40 42 41
rect 58 40 66 41
rect 82 40 90 41
rect 106 40 114 41
rect 130 40 138 41
rect 154 40 162 41
rect 178 40 186 41
rect 202 40 210 41
rect 226 40 234 41
rect 250 40 258 41
<< labels >>
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 13 44 13 44 1 GND
rlabel metal2 40 96 40 96 1 D
port 1 n
rlabel metal2 280 122 280 122 1 Q
port 4 n
rlabel metal2 264 109 264 109 1 QN
port 5 n
rlabel metal2 185 96 185 96 1 CLKN
port 6 n
<< end >>
