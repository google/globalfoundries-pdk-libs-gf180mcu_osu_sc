magic
tech gf180mcuC
timestamp 1661524996
<< nwell >>
rect 0 100 280 162
<< nmos >>
rect 19 58 25 75
rect 36 58 42 75
rect 53 58 59 75
rect 70 58 76 75
rect 87 58 93 75
rect 104 58 110 75
rect 121 58 127 75
rect 138 58 144 75
rect 155 58 161 75
rect 172 58 178 75
rect 189 58 195 75
rect 206 58 212 75
rect 223 58 229 75
rect 255 58 261 75
<< pmos >>
rect 19 109 25 143
rect 36 109 42 143
rect 53 109 59 143
rect 70 109 76 143
rect 87 109 93 143
rect 104 109 110 143
rect 121 109 127 143
rect 138 109 144 143
rect 155 109 161 143
rect 172 109 178 143
rect 189 109 195 143
rect 206 109 212 143
rect 223 109 229 143
rect 255 109 261 143
<< ndiff >>
rect 9 65 19 75
rect 9 60 11 65
rect 16 60 19 65
rect 9 58 19 60
rect 25 65 36 75
rect 25 60 28 65
rect 33 60 36 65
rect 25 58 36 60
rect 42 65 53 75
rect 42 60 45 65
rect 50 60 53 65
rect 42 58 53 60
rect 59 65 70 75
rect 59 60 62 65
rect 67 60 70 65
rect 59 58 70 60
rect 76 58 87 75
rect 93 65 104 75
rect 93 60 96 65
rect 101 60 104 65
rect 93 58 104 60
rect 110 65 121 75
rect 110 60 113 65
rect 118 60 121 65
rect 110 58 121 60
rect 127 65 138 75
rect 127 60 130 65
rect 135 60 138 65
rect 127 58 138 60
rect 144 65 155 75
rect 144 60 147 65
rect 152 60 155 65
rect 144 58 155 60
rect 161 65 172 75
rect 161 60 164 65
rect 169 60 172 65
rect 161 58 172 60
rect 178 58 189 75
rect 195 58 206 75
rect 212 65 223 75
rect 212 60 215 65
rect 220 60 223 65
rect 212 58 223 60
rect 229 65 239 75
rect 229 60 232 65
rect 237 60 239 65
rect 229 58 239 60
rect 245 65 255 75
rect 245 60 247 65
rect 252 60 255 65
rect 245 58 255 60
rect 261 65 271 75
rect 261 60 264 65
rect 269 60 271 65
rect 261 58 271 60
<< pdiff >>
rect 9 141 19 143
rect 9 135 11 141
rect 16 135 19 141
rect 9 109 19 135
rect 25 141 36 143
rect 25 135 28 141
rect 33 135 36 141
rect 25 109 36 135
rect 42 141 53 143
rect 42 135 45 141
rect 50 135 53 141
rect 42 109 53 135
rect 59 141 70 143
rect 59 136 62 141
rect 67 136 70 141
rect 59 109 70 136
rect 76 109 87 143
rect 93 141 104 143
rect 93 135 96 141
rect 101 135 104 141
rect 93 109 104 135
rect 110 141 121 143
rect 110 135 113 141
rect 118 135 121 141
rect 110 109 121 135
rect 127 141 138 143
rect 127 135 130 141
rect 135 135 138 141
rect 127 109 138 135
rect 144 141 155 143
rect 144 135 147 141
rect 152 135 155 141
rect 144 109 155 135
rect 161 128 172 143
rect 161 122 164 128
rect 169 122 172 128
rect 161 109 172 122
rect 178 109 189 143
rect 195 109 206 143
rect 212 141 223 143
rect 212 135 215 141
rect 220 135 223 141
rect 212 109 223 135
rect 229 141 239 143
rect 229 135 232 141
rect 237 135 239 141
rect 229 109 239 135
rect 245 141 255 143
rect 245 135 247 141
rect 252 135 255 141
rect 245 109 255 135
rect 261 141 271 143
rect 261 135 264 141
rect 269 135 271 141
rect 261 109 271 135
<< ndiffc >>
rect 11 60 16 65
rect 28 60 33 65
rect 45 60 50 65
rect 62 60 67 65
rect 96 60 101 65
rect 113 60 118 65
rect 130 60 135 65
rect 147 60 152 65
rect 164 60 169 65
rect 215 60 220 65
rect 232 60 237 65
rect 247 60 252 65
rect 264 60 269 65
<< pdiffc >>
rect 11 135 16 141
rect 28 135 33 141
rect 45 135 50 141
rect 62 136 67 141
rect 96 135 101 141
rect 113 135 118 141
rect 130 135 135 141
rect 147 135 152 141
rect 164 122 169 128
rect 215 135 220 141
rect 232 135 237 141
rect 247 135 252 141
rect 264 135 269 141
<< psubdiff >>
rect 9 49 18 51
rect 9 44 11 49
rect 16 44 18 49
rect 9 42 18 44
rect 33 49 42 51
rect 33 44 35 49
rect 40 44 42 49
rect 33 42 42 44
rect 57 49 66 51
rect 57 44 59 49
rect 64 44 66 49
rect 57 42 66 44
rect 81 49 90 51
rect 81 44 83 49
rect 88 44 90 49
rect 81 42 90 44
rect 105 49 114 51
rect 105 44 107 49
rect 112 44 114 49
rect 105 42 114 44
rect 129 49 138 51
rect 129 44 131 49
rect 136 44 138 49
rect 129 42 138 44
rect 153 49 162 51
rect 153 44 155 49
rect 160 44 162 49
rect 153 42 162 44
rect 177 49 186 51
rect 177 44 179 49
rect 184 44 186 49
rect 177 42 186 44
rect 201 49 210 51
rect 201 44 203 49
rect 208 44 210 49
rect 201 42 210 44
rect 225 49 234 51
rect 225 44 227 49
rect 232 44 234 49
rect 225 42 234 44
rect 249 49 258 51
rect 249 44 251 49
rect 256 44 258 49
rect 249 42 258 44
<< nsubdiff >>
rect 9 157 18 159
rect 9 152 11 157
rect 16 152 18 157
rect 9 150 18 152
rect 33 157 42 159
rect 33 152 35 157
rect 40 152 42 157
rect 33 150 42 152
rect 57 157 66 159
rect 57 152 59 157
rect 64 152 66 157
rect 57 150 66 152
rect 81 157 90 159
rect 81 152 83 157
rect 88 152 90 157
rect 81 150 90 152
rect 105 157 114 159
rect 105 152 107 157
rect 112 152 114 157
rect 105 150 114 152
rect 129 157 138 159
rect 129 152 131 157
rect 136 152 138 157
rect 129 150 138 152
rect 153 157 162 159
rect 153 152 155 157
rect 160 152 162 157
rect 153 150 162 152
rect 177 157 186 159
rect 177 152 179 157
rect 184 152 186 157
rect 177 150 186 152
rect 201 157 210 159
rect 201 152 203 157
rect 208 152 210 157
rect 201 150 210 152
rect 225 157 234 159
rect 225 152 227 157
rect 232 152 234 157
rect 225 150 234 152
rect 249 157 258 159
rect 249 152 251 157
rect 256 152 258 157
rect 249 150 258 152
<< psubdiffcont >>
rect 11 44 16 49
rect 35 44 40 49
rect 59 44 64 49
rect 83 44 88 49
rect 107 44 112 49
rect 131 44 136 49
rect 155 44 160 49
rect 179 44 184 49
rect 203 44 208 49
rect 227 44 232 49
rect 251 44 256 49
<< nsubdiffcont >>
rect 11 152 16 157
rect 35 152 40 157
rect 59 152 64 157
rect 83 152 88 157
rect 107 152 112 157
rect 131 152 136 157
rect 155 152 160 157
rect 179 152 184 157
rect 203 152 208 157
rect 227 152 232 157
rect 251 152 256 157
<< polysilicon >>
rect 19 143 25 148
rect 36 143 42 148
rect 53 143 59 148
rect 70 143 76 148
rect 87 143 93 148
rect 104 143 110 148
rect 121 143 127 148
rect 138 143 144 148
rect 155 143 161 148
rect 172 143 178 148
rect 189 143 195 148
rect 206 143 212 148
rect 223 143 229 148
rect 255 143 261 148
rect 19 91 25 109
rect 36 104 42 109
rect 30 102 42 104
rect 30 96 32 102
rect 38 96 42 102
rect 30 94 42 96
rect 12 89 25 91
rect 12 83 14 89
rect 20 83 25 89
rect 12 81 25 83
rect 19 75 25 81
rect 36 75 42 94
rect 53 91 59 109
rect 70 107 76 109
rect 87 107 93 109
rect 104 107 110 109
rect 121 107 127 109
rect 70 105 82 107
rect 70 99 74 105
rect 80 99 82 105
rect 70 97 82 99
rect 87 102 110 107
rect 115 105 127 107
rect 51 89 61 91
rect 51 83 53 89
rect 59 83 61 89
rect 51 81 61 83
rect 53 75 59 81
rect 70 75 76 97
rect 87 94 93 102
rect 115 99 117 105
rect 123 99 127 105
rect 115 97 127 99
rect 87 92 102 94
rect 87 86 94 92
rect 100 86 102 92
rect 87 84 102 86
rect 87 79 110 84
rect 87 75 93 79
rect 104 75 110 79
rect 121 75 127 97
rect 138 94 144 109
rect 155 94 161 109
rect 172 94 178 109
rect 189 107 195 109
rect 189 105 201 107
rect 189 99 193 105
rect 199 99 201 105
rect 189 97 201 99
rect 138 92 149 94
rect 138 86 141 92
rect 147 86 149 92
rect 138 84 149 86
rect 155 92 166 94
rect 155 86 158 92
rect 164 86 166 92
rect 155 84 166 86
rect 172 92 184 94
rect 172 86 176 92
rect 182 86 184 92
rect 172 84 184 86
rect 138 75 144 84
rect 155 75 161 84
rect 172 75 178 84
rect 189 75 195 97
rect 206 92 212 109
rect 223 94 229 109
rect 255 94 261 109
rect 202 90 212 92
rect 202 84 204 90
rect 210 84 212 90
rect 217 92 229 94
rect 217 86 219 92
rect 225 86 229 92
rect 217 84 229 86
rect 249 92 261 94
rect 249 86 251 92
rect 257 86 261 92
rect 249 84 261 86
rect 202 82 212 84
rect 206 75 212 82
rect 223 75 229 84
rect 255 75 261 84
rect 19 53 25 58
rect 36 53 42 58
rect 53 53 59 58
rect 70 53 76 58
rect 87 53 93 58
rect 104 53 110 58
rect 121 53 127 58
rect 138 53 144 58
rect 155 53 161 58
rect 172 53 178 58
rect 189 53 195 58
rect 206 53 212 58
rect 223 53 229 58
rect 255 53 261 58
<< polycontact >>
rect 32 96 38 102
rect 14 83 20 89
rect 74 99 80 105
rect 53 83 59 89
rect 117 99 123 105
rect 94 86 100 92
rect 193 99 199 105
rect 141 86 147 92
rect 158 86 164 92
rect 176 86 182 92
rect 204 84 210 90
rect 219 86 225 92
rect 251 86 257 92
<< metal1 >>
rect 0 157 280 162
rect 0 151 11 157
rect 17 151 35 157
rect 41 151 59 157
rect 65 151 83 157
rect 89 151 107 157
rect 113 151 131 157
rect 137 151 155 157
rect 161 151 179 157
rect 185 151 203 157
rect 209 151 227 157
rect 233 151 251 157
rect 257 151 280 157
rect 0 150 280 151
rect 11 141 16 143
rect 11 128 16 135
rect 28 141 33 150
rect 28 133 33 135
rect 45 141 50 143
rect 45 128 50 135
rect 62 141 68 143
rect 62 133 68 135
rect 96 141 101 150
rect 96 133 101 135
rect 113 141 118 143
rect 11 123 50 128
rect 113 128 118 135
rect 130 141 135 150
rect 130 133 135 135
rect 147 141 152 143
rect 147 128 152 135
rect 215 141 220 150
rect 215 133 220 135
rect 232 141 237 143
rect 113 123 152 128
rect 162 122 164 128
rect 170 122 172 128
rect 32 112 80 118
rect 32 102 38 112
rect 32 94 38 96
rect 43 101 69 107
rect 43 89 48 101
rect 64 92 69 101
rect 74 105 80 112
rect 117 111 199 117
rect 117 105 123 111
rect 80 99 117 105
rect 74 97 80 99
rect 117 97 123 99
rect 128 100 182 106
rect 128 92 134 100
rect 12 83 14 89
rect 20 83 48 89
rect 53 89 59 91
rect 64 86 94 92
rect 100 86 134 92
rect 141 92 147 94
rect 176 92 182 100
rect 193 105 199 111
rect 193 97 199 99
rect 232 106 237 135
rect 247 141 252 150
rect 247 133 252 135
rect 264 141 269 143
rect 264 106 269 135
rect 232 105 238 106
rect 264 105 273 106
rect 232 99 233 105
rect 239 99 241 105
rect 264 99 267 105
rect 273 99 275 105
rect 232 98 238 99
rect 264 98 273 99
rect 156 86 158 92
rect 164 86 166 92
rect 174 86 176 92
rect 182 86 184 92
rect 53 81 59 83
rect 141 81 147 86
rect 195 84 204 90
rect 210 84 212 90
rect 217 86 219 92
rect 225 86 227 92
rect 195 81 201 84
rect 53 75 201 81
rect 10 66 16 68
rect 10 58 16 60
rect 28 65 33 67
rect 28 51 33 60
rect 44 66 50 68
rect 44 58 50 60
rect 62 66 68 68
rect 62 58 68 60
rect 96 65 101 67
rect 96 51 101 60
rect 113 66 119 68
rect 113 58 119 60
rect 130 65 135 67
rect 130 51 135 60
rect 146 66 152 68
rect 146 58 152 60
rect 164 66 170 68
rect 164 58 170 60
rect 215 65 220 67
rect 215 51 220 60
rect 232 65 237 98
rect 249 86 251 92
rect 257 86 259 92
rect 232 58 237 60
rect 247 65 252 67
rect 247 51 252 60
rect 264 65 269 98
rect 264 58 269 60
rect 0 50 280 51
rect 0 44 11 50
rect 17 44 35 50
rect 41 44 59 50
rect 65 44 83 50
rect 89 44 107 50
rect 113 44 131 50
rect 137 44 155 50
rect 161 44 179 50
rect 185 44 203 50
rect 209 44 227 50
rect 233 44 251 50
rect 257 44 280 50
rect 0 39 280 44
<< via1 >>
rect 11 152 16 157
rect 16 152 17 157
rect 11 151 17 152
rect 35 152 40 157
rect 40 152 41 157
rect 35 151 41 152
rect 59 152 64 157
rect 64 152 65 157
rect 59 151 65 152
rect 83 152 88 157
rect 88 152 89 157
rect 83 151 89 152
rect 107 152 112 157
rect 112 152 113 157
rect 107 151 113 152
rect 131 152 136 157
rect 136 152 137 157
rect 131 151 137 152
rect 155 152 160 157
rect 160 152 161 157
rect 155 151 161 152
rect 179 152 184 157
rect 184 152 185 157
rect 179 151 185 152
rect 203 152 208 157
rect 208 152 209 157
rect 203 151 209 152
rect 227 152 232 157
rect 232 152 233 157
rect 227 151 233 152
rect 251 152 256 157
rect 256 152 257 157
rect 251 151 257 152
rect 62 136 67 141
rect 67 136 68 141
rect 62 135 68 136
rect 164 122 169 128
rect 169 122 170 128
rect 32 96 38 102
rect 14 83 20 89
rect 53 83 59 89
rect 233 99 239 105
rect 267 99 273 105
rect 158 86 164 92
rect 219 86 225 92
rect 10 65 16 66
rect 10 60 11 65
rect 11 60 16 65
rect 44 65 50 66
rect 44 60 45 65
rect 45 60 50 65
rect 62 65 68 66
rect 62 60 67 65
rect 67 60 68 65
rect 113 65 119 66
rect 113 60 118 65
rect 118 60 119 65
rect 146 65 152 66
rect 146 60 147 65
rect 147 60 152 65
rect 164 65 170 66
rect 164 60 169 65
rect 169 60 170 65
rect 251 86 257 92
rect 11 49 17 50
rect 11 44 16 49
rect 16 44 17 49
rect 35 49 41 50
rect 35 44 40 49
rect 40 44 41 49
rect 59 49 65 50
rect 59 44 64 49
rect 64 44 65 49
rect 83 49 89 50
rect 83 44 88 49
rect 88 44 89 49
rect 107 49 113 50
rect 107 44 112 49
rect 112 44 113 49
rect 131 49 137 50
rect 131 44 136 49
rect 136 44 137 49
rect 155 49 161 50
rect 155 44 160 49
rect 160 44 161 49
rect 179 49 185 50
rect 179 44 184 49
rect 184 44 185 49
rect 203 49 209 50
rect 203 44 208 49
rect 208 44 209 49
rect 227 49 233 50
rect 227 44 232 49
rect 232 44 233 49
rect 251 49 257 50
rect 251 44 256 49
rect 256 44 257 49
<< metal2 >>
rect 10 157 18 158
rect 34 157 42 158
rect 58 157 66 158
rect 82 157 90 158
rect 106 157 114 158
rect 130 157 138 158
rect 154 157 162 158
rect 178 157 186 158
rect 202 157 210 158
rect 226 157 234 158
rect 250 157 258 158
rect 9 151 11 157
rect 17 151 19 157
rect 33 151 35 157
rect 41 151 43 157
rect 57 151 59 157
rect 65 151 67 157
rect 81 151 83 157
rect 89 151 91 157
rect 105 151 107 157
rect 113 151 115 157
rect 129 151 131 157
rect 137 151 139 157
rect 153 151 155 157
rect 161 151 163 157
rect 177 151 179 157
rect 185 151 187 157
rect 201 151 203 157
rect 209 151 211 157
rect 225 151 227 157
rect 233 151 235 157
rect 249 151 251 157
rect 257 151 259 157
rect 10 150 18 151
rect 34 150 42 151
rect 58 150 66 151
rect 82 150 90 151
rect 106 150 114 151
rect 130 150 138 151
rect 154 150 162 151
rect 178 150 186 151
rect 202 150 210 151
rect 226 150 234 151
rect 250 150 258 151
rect 62 142 68 143
rect 61 141 69 142
rect 60 135 62 141
rect 68 135 257 141
rect 61 134 69 135
rect 31 102 39 103
rect 30 96 32 102
rect 38 96 40 102
rect 31 95 39 96
rect 75 92 81 135
rect 163 128 171 129
rect 162 122 164 128
rect 170 122 225 128
rect 163 121 171 122
rect 157 92 165 93
rect 12 89 22 90
rect 52 89 60 90
rect 12 83 14 89
rect 20 83 22 89
rect 51 83 53 89
rect 59 83 61 89
rect 75 86 158 92
rect 164 86 166 92
rect 12 82 22 83
rect 52 82 60 83
rect 10 67 16 68
rect 44 67 50 68
rect 62 67 68 68
rect 9 66 17 67
rect 43 66 51 67
rect 9 60 10 66
rect 16 60 44 66
rect 50 60 51 66
rect 9 59 17 60
rect 43 59 51 60
rect 61 66 69 67
rect 75 66 81 86
rect 157 85 165 86
rect 113 67 119 68
rect 146 67 152 68
rect 61 60 62 66
rect 68 60 81 66
rect 112 66 120 67
rect 145 66 153 67
rect 163 66 171 67
rect 177 66 183 122
rect 219 93 225 122
rect 232 105 240 106
rect 231 99 233 105
rect 239 99 241 105
rect 232 98 240 99
rect 251 93 257 135
rect 266 105 274 106
rect 265 99 267 105
rect 273 99 275 105
rect 266 98 274 99
rect 218 92 226 93
rect 250 92 258 93
rect 218 86 219 92
rect 225 86 226 92
rect 249 86 251 92
rect 257 86 259 92
rect 218 85 226 86
rect 250 85 258 86
rect 219 84 225 85
rect 251 84 257 85
rect 112 60 113 66
rect 119 60 146 66
rect 152 60 153 66
rect 162 60 164 66
rect 170 60 183 66
rect 61 59 69 60
rect 112 59 120 60
rect 145 59 153 60
rect 163 59 171 60
rect 10 58 16 59
rect 44 58 50 59
rect 62 58 68 59
rect 113 58 119 59
rect 146 58 152 59
rect 10 50 18 51
rect 34 50 42 51
rect 58 50 66 51
rect 82 50 90 51
rect 106 50 114 51
rect 130 50 138 51
rect 154 50 162 51
rect 178 50 186 51
rect 202 50 210 51
rect 226 50 234 51
rect 250 50 258 51
rect 9 44 11 50
rect 17 44 19 50
rect 33 44 35 50
rect 41 44 43 50
rect 57 44 59 50
rect 65 44 67 50
rect 81 44 83 50
rect 89 44 91 50
rect 105 44 107 50
rect 113 44 115 50
rect 129 44 131 50
rect 137 44 139 50
rect 153 44 155 50
rect 161 44 163 50
rect 177 44 179 50
rect 185 44 187 50
rect 201 44 203 50
rect 209 44 211 50
rect 225 44 227 50
rect 233 44 235 50
rect 249 44 251 50
rect 257 44 259 50
rect 10 43 18 44
rect 34 43 42 44
rect 58 43 66 44
rect 82 43 90 44
rect 106 43 114 44
rect 130 43 138 44
rect 154 43 162 44
rect 178 43 186 44
rect 202 43 210 44
rect 226 43 234 44
rect 250 43 258 44
<< labels >>
rlabel metal2 14 154 14 154 1 VDD
rlabel metal2 14 47 14 47 1 GND
rlabel metal2 17 86 17 86 1 A
port 7 n
rlabel metal2 35 99 35 99 1 B
port 8 n
rlabel metal2 56 86 56 86 1 CI
port 9 n
rlabel metal2 236 102 236 102 1 S
port 10 n
rlabel metal2 270 102 270 102 1 CO
port 11 n
<< end >>
