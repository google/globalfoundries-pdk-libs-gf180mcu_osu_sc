# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__xor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__xor2_1 0 0 ;
  SIZE 6.2 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 6.2 8.1 ;
        RECT 4.5 5.45 4.75 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.2 0.6 ;
        RECT 4.5 0 4.75 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.25 2.2 1.75 2.5 ;
      LAYER MET2 ;
        RECT 1.25 2.2 1.75 2.5 ;
        RECT 1.3 2.15 1.7 2.55 ;
      LAYER VIA12 ;
        RECT 1.37 2.22 1.63 2.48 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.95 3.5 5.1 3.8 ;
      LAYER MET2 ;
        RECT 4.6 3.5 5.1 3.8 ;
        RECT 4.65 3.45 5.05 3.85 ;
        RECT 1.95 3.5 2.45 3.8 ;
        RECT 2 3.45 2.4 3.85 ;
      LAYER VIA12 ;
        RECT 2.07 3.52 2.33 3.78 ;
        RECT 4.72 3.52 4.98 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.9 1.4 3.2 1.95 ;
        RECT 2.95 0.95 3.2 1.95 ;
        RECT 2.95 5.35 3.2 7.15 ;
        RECT 2.9 5.35 3.2 5.85 ;
      LAYER MET2 ;
        RECT 2.8 1.5 3.3 1.9 ;
        RECT 2.85 5.4 3.25 5.8 ;
        RECT 2.9 1.5 3.2 5.95 ;
      LAYER VIA12 ;
        RECT 2.92 5.47 3.18 5.73 ;
        RECT 2.92 1.57 3.18 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.35 0.95 5.6 7.15 ;
      RECT 2.55 4.8 5.6 5.1 ;
      RECT 4.05 2.2 5.6 2.5 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 4.15 4.05 4.45 ;
  END
END gf180mcu_osu_sc_gp12t3v3__xor2_1
