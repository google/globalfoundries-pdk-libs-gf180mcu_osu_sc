# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_oai21_1 0 0 ;
  SIZE 4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4 6.15 ;
        RECT 3.05 4.45 3.3 6.15 ;
        RECT 0.65 3.5 0.9 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4 0.6 ;
        RECT 1.35 0 1.6 1.4 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.65 2.85 2.15 3.15 ;
      LAYER MET2 ;
        RECT 1.65 2.8 2.15 3.2 ;
      LAYER VIA12 ;
        RECT 1.77 2.87 2.03 3.13 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.35 2.2 2.85 2.5 ;
      LAYER MET2 ;
        RECT 2.35 2.15 2.85 2.55 ;
      LAYER VIA12 ;
        RECT 2.47 2.22 2.73 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 3.5 3.5 3.8 ;
        RECT 3.1 3.45 3.45 3.8 ;
        RECT 3.15 0.95 3.4 3.8 ;
        RECT 2.1 3.5 2.45 5.2 ;
      LAYER MET2 ;
        RECT 3 3.5 3.5 3.8 ;
        RECT 3.05 3.45 3.45 3.85 ;
      LAYER VIA12 ;
        RECT 3.12 3.52 3.38 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.65 2.55 1.9 ;
      RECT 2.2 0.95 2.55 1.9 ;
      RECT 0.5 0.95 0.75 1.9 ;
  END
END gf180mcu_osu_sc_9T_oai21_1
