# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__dffs_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__dffs_1 0 0 ;
  SIZE 15.45 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 15.45 8.3 ;
        RECT 13.8 5.55 14.05 8.3 ;
        RECT 11.35 6.8 11.6 8.3 ;
        RECT 8.9 6.3 9.15 8.3 ;
        RECT 6.1 5.55 6.35 8.3 ;
        RECT 3.05 5.55 3.3 8.3 ;
        RECT 1.45 6.3 1.7 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 15.45 0.7 ;
        RECT 13.8 0 14.05 1.9 ;
        RECT 10.65 0 10.9 1.9 ;
        RECT 8.9 0 9.15 1.9 ;
        RECT 6.1 0 6.35 1.5 ;
        RECT 3.05 0 3.3 1.9 ;
        RECT 2.15 0 2.4 1.9 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal1 ;
        RECT 9.3 4.25 9.8 4.55 ;
        RECT 7.15 4.25 8.2 4.55 ;
        RECT 7.05 2.25 7.55 2.55 ;
        RECT 7.15 2.25 7.45 4.55 ;
        RECT 4.25 4.25 5.4 4.55 ;
        RECT 4.9 2.3 5.4 2.6 ;
        RECT 5 2.3 5.3 4.55 ;
      LAYER Metal2 ;
        RECT 4.9 4.25 9.8 4.55 ;
        RECT 9.35 4.2 9.75 4.6 ;
        RECT 7.7 4.2 8.2 4.6 ;
        RECT 4.9 4.2 5.35 4.6 ;
      LAYER Via1 ;
        RECT 5.02 4.27 5.28 4.53 ;
        RECT 7.82 4.27 8.08 4.53 ;
        RECT 9.42 4.27 9.68 4.53 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.55 3.6 4.05 3.9 ;
      LAYER Metal2 ;
        RECT 3.55 3.55 4.05 3.95 ;
      LAYER Via1 ;
        RECT 3.67 3.62 3.93 3.88 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 14.65 4.9 15.15 5.25 ;
        RECT 14.65 4.85 15.1 5.25 ;
        RECT 14.65 1.05 14.9 7.25 ;
      LAYER Metal2 ;
        RECT 14.65 4.9 15.15 5.2 ;
        RECT 14.7 4.85 15.1 5.25 ;
      LAYER Via1 ;
        RECT 14.77 4.92 15.03 5.18 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12.95 4.25 14.4 4.55 ;
        RECT 14.05 2.15 14.3 4.55 ;
        RECT 12.95 2.15 14.3 2.4 ;
        RECT 12.95 4.25 13.2 7.25 ;
        RECT 12.95 1.05 13.2 2.4 ;
      LAYER Metal2 ;
        RECT 13.9 4.25 14.4 4.55 ;
        RECT 13.95 4.2 14.35 4.6 ;
      LAYER Via1 ;
        RECT 14.02 4.27 14.28 4.53 ;
    END
  END QN
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 11.55 4.25 12.05 4.55 ;
        RECT 5.7 4.9 6.2 5.2 ;
        RECT 5.7 2.3 6.2 2.6 ;
        RECT 5.8 2.3 6.1 5.2 ;
        RECT 2.3 5.8 2.55 7.25 ;
        RECT 0.75 2.3 2.5 2.6 ;
        RECT 2.1 2.25 2.35 2.65 ;
        RECT 0.6 5.8 2.55 6.05 ;
        RECT 0.75 4.25 1.5 4.55 ;
        RECT 0.75 1.05 1 6.05 ;
        RECT 0.6 5.8 0.85 7.25 ;
      LAYER Metal2 ;
        RECT 11.55 4.2 12.05 4.6 ;
        RECT 1.1 5.55 11.95 5.85 ;
        RECT 11.65 4.2 11.95 5.85 ;
        RECT 1 4.2 1.5 4.6 ;
        RECT 1.1 4.2 1.4 5.85 ;
        RECT 2 2.3 6.2 2.6 ;
        RECT 5.75 2.25 6.15 2.65 ;
        RECT 2 2.25 2.5 2.65 ;
      LAYER Via1 ;
        RECT 1.12 4.27 1.38 4.53 ;
        RECT 2.12 2.32 2.38 2.58 ;
        RECT 5.82 2.32 6.08 2.58 ;
        RECT 11.67 4.27 11.93 4.53 ;
    END
  END SN
  OBS
    LAYER Metal2 ;
      RECT 13.2 2.9 13.6 3.3 ;
      RECT 12.85 2.95 13.65 3.25 ;
      RECT 10.55 2.2 11.05 2.6 ;
      RECT 10.55 1.65 10.95 2.6 ;
      RECT 7.45 1.6 7.85 2 ;
      RECT 7.4 1.65 10.95 1.95 ;
      RECT 10.6 4.85 11 5.25 ;
      RECT 8.4 4.85 8.8 5.25 ;
      RECT 8.35 4.9 11.05 5.2 ;
      RECT 9.7 2.9 10.1 3.3 ;
      RECT 7.75 2.9 8.15 3.3 ;
      RECT 7.7 2.95 10.2 3.25 ;
      RECT 8.45 3.55 8.85 3.95 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 12.25 4.85 12.75 5.25 ;
      RECT 2 3.55 2.5 3.95 ;
    LAYER Via1 ;
      RECT 13.27 2.97 13.53 3.23 ;
      RECT 12.37 4.92 12.63 5.18 ;
      RECT 10.67 2.27 10.93 2.53 ;
      RECT 10.67 4.92 10.93 5.18 ;
      RECT 9.77 2.97 10.03 3.23 ;
      RECT 8.52 3.62 8.78 3.88 ;
      RECT 8.47 4.92 8.73 5.18 ;
      RECT 7.82 2.97 8.08 3.23 ;
      RECT 7.52 1.67 7.78 1.93 ;
      RECT 2.12 3.62 2.38 3.88 ;
    LAYER Metal1 ;
      RECT 12.35 2.95 12.65 5.3 ;
      RECT 10.65 4.8 10.95 5.3 ;
      RECT 10.65 4.9 12.65 5.2 ;
      RECT 12.05 2.95 13.65 3.25 ;
      RECT 12.05 1.05 12.3 3.25 ;
      RECT 12.2 6.3 12.45 7.25 ;
      RECT 10.5 6.3 10.75 7.25 ;
      RECT 10.5 6.3 12.45 6.55 ;
      RECT 9.75 4.85 10 7.25 ;
      RECT 9.75 4.85 10.3 5.1 ;
      RECT 10.05 3.65 10.3 5.1 ;
      RECT 9.75 2.85 10.05 3.9 ;
      RECT 9.75 1.05 10 3.9 ;
      RECT 8.35 4.9 8.85 5.2 ;
      RECT 8.45 3.6 8.75 5.2 ;
      RECT 8.4 3.6 8.9 3.9 ;
      RECT 7.5 6.05 7.75 7.25 ;
      RECT 6.6 6.05 7.75 6.3 ;
      RECT 6.6 3.55 6.85 6.3 ;
      RECT 6.55 1.7 6.8 3.8 ;
      RECT 6.55 1.7 7.9 1.95 ;
      RECT 7.5 1.65 7.9 1.95 ;
      RECT 7.5 1.05 7.75 1.95 ;
      RECT 4.7 5.05 4.95 7.25 ;
      RECT 3.05 5.05 4.95 5.3 ;
      RECT 3.05 2.35 3.3 5.3 ;
      RECT 2 3.6 3.3 3.9 ;
      RECT 3.05 2.35 4.05 2.6 ;
      RECT 3.65 1.65 4.05 2.6 ;
      RECT 3.65 1.65 4.95 1.9 ;
      RECT 4.7 1.05 4.95 1.9 ;
      RECT 10.55 2.25 11.05 2.55 ;
      RECT 7.7 2.95 8.2 3.25 ;
  END
END gf180mcu_osu_sc_gp12t3v3__dffs_1
