##################################################################################
#
#           GLOBALFOUNDRIES
#
##################################################################################
#
# 180MCU Tech LEF File
# based on DRM DM-000013-01 Rev 13
# TFG-Version: 2.1.9
# Date: February 2018
#-------------------------------------------------------
# metal stack option: 5LM_1TM_9K
# Preferred routing directions:
# vertical:   MET2 MET4 
# horizontal: MET1 MET3 MET5
#------------------------------------------------------
# This Techfile contains not correct Parasitic Information.
# USE Appropriate parasitic files for Parasitic Extraction.
#------------------------------------------------------

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000  ;
    CAPACITANCE PICOFARADS 1 ;
    CURRENT MILLIAMPS 1 ;
    RESISTANCE OHMS 1 ;
END UNITS

PROPERTYDEFINITIONS
  LAYER LEF58_EOLENCLOSURE STRING ;
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

MANUFACTURINGGRID 0.0050 ;
CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS ON ;

LAYER POLY2
 TYPE MASTERSLICE ;
END POLY2

LAYER CONT
 TYPE CUT ;
END CONT


LAYER MET1
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.56 ; 
    OFFSET 0.28 ;

    MINWIDTH 0.230 ;                   # Mn.1  (n=1)
    WIDTH 0.230 ;                      # Mn.1  (n=1)
    SPACING 0.230  ;                   # Mn.2a (n=1)
    SPACING 0.300 RANGE 10.005 999.00 ; # Mn.2b
    AREA 0.1444 ;                      # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNASIDEAREARATIO 400 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END MET1


LAYER VIA12
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.00 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;
  PROPERTY LEF58_EOLENCLOSURE "
  	EOLENCLOSURE 0.34 0.06 ;" ; 

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END VIA12


LAYER MET2
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.56 ; 
    OFFSET 0.28 ;

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END MET2


LAYER VIA23
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END VIA23


LAYER MET3
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    PITCH 0.56 ; 
    OFFSET 0.28 ;

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END MET3


LAYER VIA34
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END VIA34


LAYER MET4
    TYPE ROUTING ;
    DIRECTION VERTICAL ;

    PITCH 0.56 ; 
    OFFSET 0.28 ;

    MINWIDTH 0.280 ;
    WIDTH 0.280 ;                        # Mn.1  (n>1)
    SPACING 0.280 ;                      # Mn.2a (n>1)
    SPACING 0.300 RANGE 10.005 999.00 ;  # Mn.2b
    AREA 0.1444 ;                        # Mn.3

    THICKNESS 0.54 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    DCCURRENTDENSITY AVERAGE 0.67 ;
    ACCURRENTDENSITY AVERAGE 1.00 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;
    RESISTANCE RPERSQ 0.090000 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END MET4


LAYER VIA45
  TYPE CUT ;
  SPACING 0.26 ;
  WIDTH   0.26 ;

  ENCLOSURE BELOW 0.01 0.06 ;
 # ENCLOSURE ABOVE 0.01 0.09 ;
  ENCLOSURE ABOVE 0.01 0.06 ;

  # a bit conservative for Vn.3/4a without considering the protrusion length of 0.28
  PROPERTY LEF58_EOLENCLOSURE " EOLENCLOSURE 0.34 0.06 ; " ;

  ARRAYSPACING CUTSPACING 0.36 ARRAYCUTS 4 SPACING 0.36 ; # Vn.2b

  ACCURRENTDENSITY AVERAGE 0.28 ;
  DCCURRENTDENSITY AVERAGE 0.18 ;
  ANTENNAMODEL OXIDE1 ;
  ANTENNAAREARATIO 20.0 ;
END VIA45



LAYER MET5
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;

    OFFSET 0.45 ;


    PITCH 0.9 ;
    MINWIDTH 0.440 ;
    WIDTH   0.440 ;                      # MT.1
    AREA    0.5625 ;                     # MT.4
    SPACING 0.460 ;                      # MT.2a
    SPACING 0.600 RANGE 10.005 999.00 ;  # MT.2b

    DCCURRENTDENSITY AVERAGE 1.21 ;
    ACCURRENTDENSITY AVERAGE 1.82 ;
    RESISTANCE RPERSQ 0.04000 ;

    THICKNESS 0.99 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO 400 ;
    ANTENNAGATEPLUSDIFF 2 ;

    CAPACITANCE CPERSQDIST 0.0000394 ;

    MINIMUMDENSITY 30.0 ;
    DENSITYCHECKWINDOW 200.0 200.0 ;
    DENSITYCHECKSTEP 100.0 ;

END MET5



LAYER OverlapCheck
 TYPE OVERLAP ;
END OverlapCheck
LAYER OBS
 TYPE MASTERSLICE ;
END OBS

LAYER PR_bndry
    TYPE MASTERSLICE ;
END PR_bndry

#------------------------------------------------------------
#  CONT VIA SECTION 
#------------------------------------------------------------
#VIA CONT1 DEFAULT
# RESISTANCE 13.5 ;
# LAYER CONT ;
# RECT -0.11 -0.11 0.11 0.11 ;
# LAYER POLY2 ;
# RECT -0.18 -0.18 0.18 0.18 ;
# LAYER MET1 ;
# RECT -0.115 -0.115 0.115 0.115 ;
#END CONT1

#VIARULE CONT1 GENERATE
# LAYER POLY2 ;
# DIRECTION HORIZONTAL ;
# OVERHANG 0.07 ;
# LAYER MET1 ;
# DIRECTION VERTICAL ;
# OVERHANG 0.005 ;
# LAYER CONT ;
# RECT -0.11 -0.11 0.11 0.11 ;
# SPACING 0.47 BY 0.47 ;
# RESISTANCE 13.5 ;
#END CONT1



#------------------------------------------------------------
#  VIA12 VIA SECTION 
#------------------------------------------------------------
 VIA VIA12_HH  DEFAULT
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER MET2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA12_HH 
 
 VIA VIA12_HV  DEFAULT
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA12_HV 
 
 VIA VIA12_VH  DEFAULT
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER MET2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA12_VH 
 
 VIA VIA12_VV  DEFAULT
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.130 -0.190 0.130 0.190 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA12_VV 
 
 VIA V12A  DEFAULT
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER MET2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END V12A 
 
 VIA V12B 
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.190 -0.130 0.190 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END V12B 
 
 VIA V12_fat 
 LAYER VIA12 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET1 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 LAYER MET2 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 RESISTANCE 5.000 ;
 END V12_fat 
 
 VIA VIA12_2CUT_H
 LAYER VIA12 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER MET1 ;
 RECT -0.450 -0.130 0.450 0.130 ;
 LAYER MET2 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 END VIA12_2CUT_H
 
 VIA VIA12_2CUT_V
 LAYER VIA12 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER MET1 ;
 RECT -0.190 -0.390 0.190 0.390 ;
 LAYER MET2 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 END VIA12_2CUT_V
 
 VIA VIA12_2X2_0_60_10_60_H_H  DEFAULT
 LAYER VIA12 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER MET2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA12_2X2_0_60_10_60_H_H 
 
 VIA VIA12_2X2_0_60_10_60_H_V  DEFAULT
 LAYER VIA12 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET1 ;
 RECT -0.450 -0.390 0.450 0.390 ;
 LAYER MET2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA12_2X2_0_60_10_60_H_V 
 
 VIA VIA12_2X2_0_60_10_60_V_H  DEFAULT
 LAYER VIA12 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER MET2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA12_2X2_0_60_10_60_V_H 
 
 VIA VIA12_2X2_0_60_10_60_V_V  DEFAULT
 LAYER VIA12 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET1 ;
 RECT -0.390 -0.450 0.390 0.450 ;
 LAYER MET2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA12_2X2_0_60_10_60_V_V 
 
VIARULE VIA12_GEN_HH GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER MET2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA12_GEN_HH

VIARULE VIA12_GEN_HV GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.060 0.000 ;
  LAYER MET2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA12_GEN_HV

VIARULE VIA12_GEN_VH GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER MET2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA12_GEN_VH

VIARULE VIA12_GEN_VV GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.000 0.060 ;
  LAYER MET2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA12_GEN_VV

VIARULE V12B GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET2 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V12B

VIARULE V12_fat GENERATE
  LAYER MET1 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET2 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA12 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V12_fat

 VIA VIA12_4X4H_HH_DEFAULT  DEFAULT
 LAYER VIA12 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER MET2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA12_4X4H_HH_DEFAULT 
 
 VIA VIA12_4X4H_HV_DEFAULT  DEFAULT
 LAYER VIA12 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET1 ;
 RECT -1.120 -1.060 1.120 1.060 ;
 LAYER MET2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA12_4X4H_HV_DEFAULT 
 
 VIA VIA12_4X4H_VH_DEFAULT  DEFAULT
 LAYER VIA12 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER MET2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA12_4X4H_VH_DEFAULT 
 
 VIA VIA12_4X4H_VV_DEFAULT  DEFAULT
 LAYER VIA12 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET1 ;
 RECT -1.060 -1.120 1.060 1.120 ;
 LAYER MET2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA12_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  VIA23 VIA SECTION 
#------------------------------------------------------------
 VIA VIA23_HH  DEFAULT
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA23_HH 
 
 VIA VIA23_HV  DEFAULT
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA23_HV 
 
 VIA VIA23_VH  DEFAULT
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA23_VH 
 
 VIA VIA23_VV  DEFAULT
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA23_VV 
 
 VIA V23B  DEFAULT
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END V23B 
 
 VIA V23A 
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END V23A 
 
 VIA V23_fat 
 LAYER VIA23 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET2 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 LAYER MET3 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 RESISTANCE 5.000 ;
 END V23_fat 
 
 VIA VIA23_2CUT_H
 LAYER VIA23 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER MET2 ;
 RECT -0.390 -0.190 0.390 0.190 ;
 LAYER MET3 ;
 RECT -0.450 -0.140 0.450 0.140 ;
 END VIA23_2CUT_H
 
 VIA VIA23_2CUT_V
 LAYER VIA23 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER MET2 ;
 RECT -0.130 -0.450 0.130 0.450 ;
 LAYER MET3 ;
 RECT -0.190 -0.400 0.190 0.400 ;
 END VIA23_2CUT_V
 
 VIA VIA23_2X2_10_60_10_60_H_H  DEFAULT
 LAYER VIA23 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA23_2X2_10_60_10_60_H_H 
 
 VIA VIA23_2X2_10_60_10_60_H_V  DEFAULT
 LAYER VIA23 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET2 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA23_2X2_10_60_10_60_H_V 
 
 VIA VIA23_2X2_10_60_10_60_V_H  DEFAULT
 LAYER VIA23 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA23_2X2_10_60_10_60_V_H 
 
 VIA VIA23_2X2_10_60_10_60_V_V  DEFAULT
 LAYER VIA23 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET2 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA23_2X2_10_60_10_60_V_V 
 
VIARULE VIA23_GEN_HH GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA23_GEN_HH

VIARULE VIA23_GEN_HV GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA23_GEN_HV

VIARULE VIA23_GEN_VH GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA23_GEN_VH

VIARULE VIA23_GEN_VV GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA23_GEN_VV

VIARULE V23B GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET3 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V23B

VIARULE V23_fat GENERATE
  LAYER MET2 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET3 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA23 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V23_fat

 VIA VIA23_4X4H_HH_DEFAULT  DEFAULT
 LAYER VIA23 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA23_4X4H_HH_DEFAULT 
 
 VIA VIA23_4X4H_HV_DEFAULT  DEFAULT
 LAYER VIA23 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET2 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA23_4X4H_HV_DEFAULT 
 
 VIA VIA23_4X4H_VH_DEFAULT  DEFAULT
 LAYER VIA23 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA23_4X4H_VH_DEFAULT 
 
 VIA VIA23_4X4H_VV_DEFAULT  DEFAULT
 LAYER VIA23 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET2 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA23_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  VIA34 VIA SECTION 
#------------------------------------------------------------
 VIA VIA34_HH  DEFAULT
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA34_HH 
 
 VIA VIA34_HV  DEFAULT
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA34_HV 
 
 VIA VIA34_VH  DEFAULT
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA34_VH 
 
 VIA VIA34_VV  DEFAULT
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA34_VV 
 
 VIA V34A  DEFAULT
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END V34A 
 
 VIA V34B 
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END V34B 
 
 VIA V34_fat 
 LAYER VIA34 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET3 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 LAYER MET4 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 RESISTANCE 5.000 ;
 END V34_fat 
 
 VIA VIA34_2CUT_H
 LAYER VIA34 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER MET3 ;
 RECT -0.450 -0.130 0.450 0.130 ;
 LAYER MET4 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 END VIA34_2CUT_H
 
 VIA VIA34_2CUT_V
 LAYER VIA34 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER MET3 ;
 RECT -0.190 -0.390 0.190 0.390 ;
 LAYER MET4 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 END VIA34_2CUT_V
 
 VIA VIA34_2X2_10_60_10_60_H_H  DEFAULT
 LAYER VIA34 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA34_2X2_10_60_10_60_H_H 
 
 VIA VIA34_2X2_10_60_10_60_H_V  DEFAULT
 LAYER VIA34 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET3 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA34_2X2_10_60_10_60_H_V 
 
 VIA VIA34_2X2_10_60_10_60_V_H  DEFAULT
 LAYER VIA34 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA34_2X2_10_60_10_60_V_H 
 
 VIA VIA34_2X2_10_60_10_60_V_V  DEFAULT
 LAYER VIA34 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET3 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA34_2X2_10_60_10_60_V_V 
 
VIARULE VIA34_GEN_HH GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA34_GEN_HH

VIARULE VIA34_GEN_HV GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA34_GEN_HV

VIARULE VIA34_GEN_VH GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA34_GEN_VH

VIARULE VIA34_GEN_VV GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA34_GEN_VV

VIARULE V34B GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET4 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V34B

VIARULE V34_fat GENERATE
  LAYER MET3 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET4 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA34 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V34_fat

 VIA VIA34_4X4H_HH_DEFAULT  DEFAULT
 LAYER VIA34 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA34_4X4H_HH_DEFAULT 
 
 VIA VIA34_4X4H_HV_DEFAULT  DEFAULT
 LAYER VIA34 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET3 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA34_4X4H_HV_DEFAULT 
 
 VIA VIA34_4X4H_VH_DEFAULT  DEFAULT
 LAYER VIA34 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA34_4X4H_VH_DEFAULT 
 
 VIA VIA34_4X4H_VV_DEFAULT  DEFAULT
 LAYER VIA34 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET3 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA34_4X4H_VV_DEFAULT 
 
#------------------------------------------------------------
#  VIA45 VIA SECTION 
#------------------------------------------------------------
 VIA VIA45_HH  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET5 ;
 RECT -0.220 -0.140 0.220 0.140 ;
 END VIA45_HH 
 
 VIA VIA45_HV  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET5 ;
 RECT -0.140 -0.220 0.140 0.220 ;
 END VIA45_HV 
 
 VIA VIA45_VH  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET5 ;
 RECT -0.220 -0.140 0.220 0.140 ;
 END VIA45_VH 
 
 VIA VIA45_VV  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET5 ;
 RECT -0.140 -0.220 0.140 0.220 ;
 END VIA45_VV 
 
 VIA V45A 
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.180 0.190 0.180 ;
 LAYER MET5 ;
 RECT -0.180 -0.190 0.180 0.190 ;
 END V45A 
 
 VIA V45B  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.180 -0.190 0.180 0.190 ;
 LAYER MET5 ;
 RECT -0.180 -0.190 0.180 0.190 ;
 END V45B 
 
 VIA VIA45_1_HH  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET5 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA45_1_HH 
 
 VIA VIA45_1_HV  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 LAYER MET5 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA45_1_HV 
 
 VIA VIA45_1_VH  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET5 ;
 RECT -0.190 -0.140 0.190 0.140 ;
 END VIA45_1_VH 
 
 VIA VIA45_1_VV  DEFAULT
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 LAYER MET5 ;
 RECT -0.140 -0.190 0.140 0.190 ;
 END VIA45_1_VV 
 
 VIA V45_fat 
 LAYER VIA45 ;
 RECT -0.130 -0.130 0.130 0.130 ;
 LAYER MET4 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 LAYER MET5 ;
 RECT -0.190 -0.190 0.190 0.190 ;
 RESISTANCE 5.000 ;
 END V45_fat 
 
 VIA VIA45_2CUT_H
 LAYER VIA45 ;
 RECT -0.390 -0.130 -0.130 0.130 ;
 RECT 0.130 -0.130 0.390 0.130 ;
 LAYER MET4 ;
 RECT -0.400 -0.190 0.400 0.190 ;
 LAYER MET5 ;
 RECT -0.450 -0.140 0.450 0.140 ;
 END VIA45_2CUT_H
 
 VIA VIA45_2CUT_V
 LAYER VIA45 ;
 RECT -0.130 -0.390 0.130 -0.130 ;
 RECT -0.130 0.130 0.130 0.390 ;
 LAYER MET4 ;
 RECT -0.140 -0.450 0.140 0.450 ;
 LAYER MET5 ;
 RECT -0.190 -0.400 0.190 0.400 ;
 END VIA45_2CUT_V
 
 VIA VIA45_2X2_10_60_10_60_H_H  DEFAULT
 LAYER VIA45 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET5 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA45_2X2_10_60_10_60_H_H 
 
 VIA VIA45_2X2_10_60_10_60_H_V  DEFAULT
 LAYER VIA45 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET4 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 LAYER MET5 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA45_2X2_10_60_10_60_H_V 
 
 VIA VIA45_2X2_10_60_10_60_V_H  DEFAULT
 LAYER VIA45 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET5 ;
 RECT -0.450 -0.400 0.450 0.400 ;
 END VIA45_2X2_10_60_10_60_V_H 
 
 VIA VIA45_2X2_10_60_10_60_V_V  DEFAULT
 LAYER VIA45 ;
 RECT -0.390 -0.390 -0.130 -0.130 ;
 RECT 0.130 -0.390 0.390 -0.130 ;
 RECT -0.390 0.130 -0.130 0.390 ;
 RECT 0.130 0.130 0.390 0.390 ;
 LAYER MET4 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 LAYER MET5 ;
 RECT -0.400 -0.450 0.400 0.450 ;
 END VIA45_2X2_10_60_10_60_V_V 
 
VIARULE VIA45_GEN_HH GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET5 ;
    ENCLOSURE 0.090 0.010 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_HH

VIARULE VIA45_GEN_HV GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET5 ;
    ENCLOSURE 0.010 0.090 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_HV

VIARULE VIA45_GEN_VH GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.090 0.010 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_VH

VIARULE VIA45_GEN_VV GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.010 0.090 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_VV

VIARULE VIA45_GEN_1_HH GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET5 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_1_HH

VIARULE VIA45_GEN_1_HV GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER MET5 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_1_HV

VIARULE VIA45_GEN_1_VH GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.060 0.010 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_1_VH

VIARULE VIA45_GEN_1_VV GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.010 0.060 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END VIA45_GEN_1_VV

VIARULE V45B GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V45B

VIARULE V45_fat GENERATE
  LAYER MET4 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER MET5 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER VIA45 ;
    RECT -0.130 -0.130 0.130 0.130 ;
    SPACING 0.520 BY 0.520 ;
END V45_fat

 VIA VIA45_4X4H_HH_DEFAULT  DEFAULT
 LAYER VIA45 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET5 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA45_4X4H_HH_DEFAULT 
 
 VIA VIA45_4X4H_HV_DEFAULT  DEFAULT
 LAYER VIA45 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET4 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 LAYER MET5 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA45_4X4H_HV_DEFAULT 
 
 VIA VIA45_4X4H_VH_DEFAULT  DEFAULT
 LAYER VIA45 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET5 ;
 RECT -1.120 -1.070 1.120 1.070 ;
 END VIA45_4X4H_VH_DEFAULT 
 
 VIA VIA45_4X4H_VV_DEFAULT  DEFAULT
 LAYER VIA45 ;
 RECT -1.060 -1.060 -0.800 -0.800 ;
 RECT -0.440 -1.060 -0.180 -0.800 ;
 RECT 0.180 -1.060 0.440 -0.800 ;
 RECT 0.800 -1.060 1.060 -0.800 ;
 RECT -1.060 -0.440 -0.800 -0.180 ;
 RECT -0.440 -0.440 -0.180 -0.180 ;
 RECT 0.180 -0.440 0.440 -0.180 ;
 RECT 0.800 -0.440 1.060 -0.180 ;
 RECT -1.060 0.180 -0.800 0.440 ;
 RECT -0.440 0.180 -0.180 0.440 ;
 RECT 0.180 0.180 0.440 0.440 ;
 RECT 0.800 0.180 1.060 0.440 ;
 RECT -1.060 0.800 -0.800 1.060 ;
 RECT -0.440 0.800 -0.180 1.060 ;
 RECT 0.180 0.800 0.440 1.060 ;
 RECT 0.800 0.800 1.060 1.060 ;
 LAYER MET4 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 LAYER MET5 ;
 RECT -1.070 -1.120 1.070 1.120 ;
 END VIA45_4X4H_VV_DEFAULT 
 

END LIBRARY
