magic
tech gf180mcuC
timestamp 1659356686
<< nwell >>
rect 0 97 77 159
<< nmos >>
rect 18 16 24 33
rect 35 16 41 33
rect 52 16 58 33
<< pmos >>
rect 21 106 27 140
rect 33 106 39 140
rect 50 106 56 140
<< ndiff >>
rect 8 25 18 33
rect 8 18 10 25
rect 15 18 18 25
rect 8 16 18 18
rect 24 25 35 33
rect 24 18 27 25
rect 32 18 35 25
rect 24 16 35 18
rect 41 25 52 33
rect 41 18 44 25
rect 49 18 52 25
rect 41 16 52 18
rect 58 31 68 33
rect 58 18 61 31
rect 66 18 68 31
rect 58 16 68 18
<< pdiff >>
rect 11 138 21 140
rect 11 108 13 138
rect 18 108 21 138
rect 11 106 21 108
rect 27 106 33 140
rect 39 138 50 140
rect 39 108 42 138
rect 47 108 50 138
rect 39 106 50 108
rect 56 138 66 140
rect 56 108 59 138
rect 64 108 66 138
rect 56 106 66 108
<< ndiffc >>
rect 10 18 15 25
rect 27 18 32 25
rect 44 18 49 25
rect 61 18 66 31
<< pdiffc >>
rect 13 108 18 138
rect 42 108 47 138
rect 59 108 64 138
<< psubdiff >>
rect 9 7 18 9
rect 9 2 11 7
rect 16 2 18 7
rect 9 0 18 2
rect 33 7 42 9
rect 33 2 35 7
rect 40 2 42 7
rect 33 0 42 2
rect 57 7 66 9
rect 57 2 59 7
rect 64 2 66 7
rect 57 0 66 2
<< nsubdiff >>
rect 9 154 18 156
rect 9 149 11 154
rect 16 149 18 154
rect 9 147 18 149
rect 33 154 42 156
rect 33 149 35 154
rect 40 149 42 154
rect 33 147 42 149
rect 57 154 66 156
rect 57 149 59 154
rect 64 149 66 154
rect 57 147 66 149
<< psubdiffcont >>
rect 11 2 16 7
rect 35 2 40 7
rect 59 2 64 7
<< nsubdiffcont >>
rect 11 149 16 154
rect 35 149 40 154
rect 59 149 64 154
<< polysilicon >>
rect 21 140 27 145
rect 33 140 39 145
rect 50 140 56 145
rect 21 104 27 106
rect 16 100 27 104
rect 16 75 22 100
rect 33 88 39 106
rect 27 86 39 88
rect 27 80 31 86
rect 37 80 39 86
rect 27 78 39 80
rect 8 73 22 75
rect 8 67 11 73
rect 17 67 22 73
rect 8 65 22 67
rect 16 42 22 65
rect 33 42 39 78
rect 50 75 56 106
rect 44 73 56 75
rect 44 67 46 73
rect 52 67 56 73
rect 44 65 56 67
rect 50 42 56 65
rect 16 39 24 42
rect 33 39 41 42
rect 50 39 58 42
rect 18 33 24 39
rect 35 33 41 39
rect 52 33 58 39
rect 18 11 24 16
rect 35 11 41 16
rect 52 11 58 16
<< polycontact >>
rect 31 80 37 86
rect 11 67 17 73
rect 46 67 52 73
<< metal1 >>
rect 0 154 77 159
rect 0 148 11 154
rect 17 148 35 154
rect 41 148 59 154
rect 65 148 77 154
rect 0 147 77 148
rect 13 138 18 147
rect 13 106 18 108
rect 42 138 47 140
rect 42 99 47 108
rect 59 138 64 147
rect 59 106 64 108
rect 42 93 59 99
rect 65 93 67 99
rect 29 80 31 86
rect 37 80 39 86
rect 9 67 11 73
rect 17 67 19 73
rect 44 67 46 73
rect 52 67 54 73
rect 59 47 64 93
rect 59 42 66 47
rect 10 32 49 37
rect 10 25 15 32
rect 10 16 15 18
rect 27 25 32 27
rect 27 9 32 18
rect 44 25 49 32
rect 44 16 49 18
rect 61 31 66 42
rect 61 16 66 18
rect 0 8 77 9
rect 0 2 11 8
rect 17 2 35 8
rect 41 2 59 8
rect 65 2 77 8
rect 0 -3 77 2
<< via1 >>
rect 11 149 16 154
rect 16 149 17 154
rect 11 148 17 149
rect 35 149 40 154
rect 40 149 41 154
rect 35 148 41 149
rect 59 149 64 154
rect 64 149 65 154
rect 59 148 65 149
rect 59 93 65 99
rect 31 80 37 86
rect 11 67 17 73
rect 46 67 52 73
rect 11 7 17 8
rect 11 2 16 7
rect 16 2 17 7
rect 35 7 41 8
rect 35 2 40 7
rect 40 2 41 7
rect 59 7 65 8
rect 59 2 64 7
rect 64 2 65 7
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 9 148 11 154
rect 17 148 19 154
rect 33 148 35 154
rect 41 148 43 154
rect 57 148 59 154
rect 65 148 67 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 57 99 67 100
rect 57 93 59 99
rect 65 93 67 99
rect 57 92 67 93
rect 29 86 39 87
rect 29 80 31 86
rect 37 80 39 86
rect 29 79 39 80
rect 9 73 19 74
rect 9 67 11 73
rect 17 67 19 73
rect 9 66 19 67
rect 44 73 54 74
rect 44 67 46 73
rect 52 67 54 73
rect 44 66 54 67
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 9 2 11 8
rect 17 2 19 8
rect 33 2 35 8
rect 41 2 43 8
rect 57 2 59 8
rect 65 2 67 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
<< labels >>
rlabel metal2 14 5 14 5 1 GND
rlabel metal2 14 151 14 151 1 VDD
rlabel metal2 34 83 34 83 1 A1
port 6 n
rlabel metal2 49 70 49 70 1 B
port 7 n
rlabel metal2 62 96 62 96 1 Y
port 4 n
rlabel metal2 14 70 14 70 1 A0
port 5 n
<< end >>
