# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__lshifup 0 0 ;
  SIZE 7.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 2.3 8.3 ;
        RECT 0.55 5.55 0.85 8.3 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal1 ;
        RECT 2.9 7.6 7.8 8.3 ;
        RECT 6.05 5.55 6.35 8.3 ;
        RECT 4.35 5.55 4.65 8.3 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 7.8 0.7 ;
        RECT 6.05 0 6.35 1.9 ;
        RECT 4.35 0 4.65 1.9 ;
        RECT 0.55 0 0.85 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 4 2.3 4.5 2.6 ;
        RECT 0.6 2.3 1.1 2.6 ;
      LAYER Metal2 ;
        RECT 4 2.25 4.5 2.65 ;
        RECT 0.6 2.3 4.5 2.6 ;
        RECT 0.6 2.25 1.1 2.65 ;
      LAYER Via1 ;
        RECT 0.72 2.32 0.98 2.58 ;
        RECT 4.12 2.32 4.38 2.58 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.9 4.25 7.3 4.55 ;
        RECT 6.95 1.05 7.25 7.25 ;
      LAYER Metal2 ;
        RECT 6.85 4.2 7.35 4.6 ;
      LAYER Via1 ;
        RECT 6.97 4.27 7.23 4.53 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 6.1 4.85 6.6 5.25 ;
      RECT 4.55 4.85 4.95 5.25 ;
      RECT 4.5 4.9 6.6 5.2 ;
      RECT 4.5 2.95 5 3.35 ;
      RECT 1.35 2.95 1.85 3.35 ;
      RECT 1.35 3 5 3.3 ;
    LAYER Via1 ;
      RECT 6.22 4.92 6.48 5.18 ;
      RECT 4.62 3.02 4.88 3.28 ;
      RECT 4.62 4.92 4.88 5.18 ;
      RECT 1.47 3.02 1.73 3.28 ;
    LAYER Metal1 ;
      RECT 5.25 1.05 5.55 7.25 ;
      RECT 4.8 4.1 5.55 4.55 ;
      RECT 3.45 1.05 3.75 7.25 ;
      RECT 4.55 4.85 5 5.3 ;
      RECT 3.45 4.9 5 5.2 ;
      RECT 1.45 1.05 1.75 7.25 ;
      RECT 1.35 3 1.85 3.3 ;
      RECT 6.1 4.9 6.6 5.2 ;
      RECT 4.5 3 5 3.3 ;
  END
END gf180mcu_osu_sc_gp12t3v3__lshifup
