magic
tech gf180mcuC
timestamp 1661875030
<< error_p >>
rect 8 61 18 123
<< nwell >>
rect 0 61 8 123
<< metal1 >>
rect 0 111 8 123
rect 0 0 8 12
<< labels >>
rlabel metal1 4 117 4 117 3 VDD
rlabel metal1 7 5 7 5 1 GND
<< end >>
