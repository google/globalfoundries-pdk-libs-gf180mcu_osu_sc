# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__xnor2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__xnor2_1 0 0 ;
  SIZE 6.4 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 6.4 6.15 ;
        RECT 4.7 4.6 4.95 6.15 ;
        RECT 1.4 4.6 1.65 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.4 0.6 ;
        RECT 4.7 0 4.95 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.5 3 4 3.3 ;
        RECT 1.25 2.2 1.75 2.5 ;
      LAYER MET2 ;
        RECT 3.55 2.95 4 3.35 ;
        RECT 3.7 0.9 4 3.35 ;
        RECT 3.6 2.9 3.95 3.4 ;
        RECT 1.35 0.9 4 1.2 ;
        RECT 1.3 2.15 1.7 2.55 ;
        RECT 1.35 0.9 1.65 2.6 ;
      LAYER VIA12 ;
        RECT 1.37 2.22 1.63 2.48 ;
        RECT 3.62 3.02 3.88 3.28 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 4.55 2.2 5.05 2.5 ;
      LAYER MET2 ;
        RECT 4.55 2.2 5.05 2.5 ;
        RECT 4.6 2.15 5 2.55 ;
        RECT 4.65 2.1 4.95 2.6 ;
      LAYER VIA12 ;
        RECT 4.67 2.22 4.93 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 1.4 3.3 1.95 ;
        RECT 3.05 0.95 3.3 1.95 ;
        RECT 3.05 4.05 3.3 5.2 ;
        RECT 3 4.05 3.3 4.75 ;
      LAYER MET2 ;
        RECT 2.9 1.5 3.4 1.9 ;
        RECT 2.95 4.1 3.35 4.5 ;
        RECT 3 4.05 3.3 4.75 ;
        RECT 2.95 1.5 3.25 4.5 ;
      LAYER VIA12 ;
        RECT 3.02 4.17 3.28 4.43 ;
        RECT 3.02 1.57 3.28 1.83 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 5.55 0.95 5.8 5.2 ;
      RECT 2.75 3.55 5.8 3.8 ;
      RECT 2.75 2.9 3.05 3.8 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 3 2.4 3.3 ;
      RECT 2.1 2.2 2.4 3.3 ;
      RECT 2.1 2.2 3.5 2.5 ;
  END
END gf180mcu_osu_sc_gp9t3v3__xnor2_1
