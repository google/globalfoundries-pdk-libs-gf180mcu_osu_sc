magic
tech gf180mcuC
timestamp 1659394415
<< nwell >>
rect 0 97 176 159
<< metal1 >>
rect 0 147 176 159
rect 0 -3 176 9
<< end >>
