* NGSPICE file created from gf180mcu_osu_sc_12T_or2_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 VDD B a_25_106# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_25_106# A a_9_106# VDD pmos_3p3 w=1.7u l=0.3u
X2 Y a_9_106# GND GND nmos_3p3 w=0.85u l=0.3u
X3 a_9_106# A GND GND nmos_3p3 w=0.85u l=0.3u
X4 Y a_9_106# VDD VDD pmos_3p3 w=1.7u l=0.3u
X5 GND B a_9_106# GND nmos_3p3 w=0.85u l=0.3u
