VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_dlatn_1
  CLASS CORE ;
  ORIGIN 7.75 0 ;
  FOREIGN gf180mcu_osu_sc_12T_dlatn_1 -7.75 0 ;
  SIZE 9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE 12T ;
  PIN CLKN
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT -2.55 4.15 -2.05 4.45 ;
        RECT -4.3 4.15 -3.8 4.45 ;
      LAYER MET2 ;
        RECT -2.55 4.1 -2.05 4.5 ;
        RECT -4.3 4.15 -2.05 4.45 ;
        RECT -4.25 4.1 -3.85 4.5 ;
      LAYER VIA12 ;
        RECT -4.18 4.17 -3.92 4.43 ;
        RECT -2.43 4.17 -2.17 4.43 ;
    END
  END CLKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -5.9 4.15 -5.4 4.45 ;
      LAYER MET2 ;
        RECT -5.9 4.1 -5.4 4.5 ;
      LAYER VIA12 ;
        RECT -5.78 4.17 -5.52 4.43 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 4.8 0.9 5.1 ;
        RECT 0.4 4.75 0.8 5.15 ;
        RECT 0.4 0.95 0.65 7.15 ;
      LAYER MET2 ;
        RECT 0.4 4.8 0.9 5.1 ;
        RECT 0.45 4.75 0.85 5.15 ;
      LAYER VIA12 ;
        RECT 0.52 4.82 0.78 5.08 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -7.75 7.5 1.25 8.1 ;
        RECT -0.45 5.45 -0.2 8.1 ;
        RECT -2.9 5.45 -2.65 8.1 ;
        RECT -6.3 6.25 -6.05 8.1 ;
      LAYER MET2 ;
        RECT -0.1 7.55 0.4 7.85 ;
        RECT -0.05 7.5 0.35 7.9 ;
        RECT -1.3 7.55 -0.8 7.85 ;
        RECT -1.25 7.5 -0.85 7.9 ;
        RECT -2.5 7.55 -2 7.85 ;
        RECT -2.45 7.5 -2.05 7.9 ;
        RECT -3.7 7.55 -3.2 7.85 ;
        RECT -3.65 7.5 -3.25 7.9 ;
        RECT -4.9 7.55 -4.4 7.85 ;
        RECT -4.85 7.5 -4.45 7.9 ;
        RECT -6.1 7.55 -5.6 7.85 ;
        RECT -6.05 7.5 -5.65 7.9 ;
        RECT -7.3 7.55 -6.8 7.85 ;
        RECT -7.25 7.5 -6.85 7.9 ;
      LAYER VIA12 ;
        RECT -7.18 7.57 -6.92 7.83 ;
        RECT -5.98 7.57 -5.72 7.83 ;
        RECT -4.78 7.57 -4.52 7.83 ;
        RECT -3.58 7.57 -3.32 7.83 ;
        RECT -2.38 7.57 -2.12 7.83 ;
        RECT -1.18 7.57 -0.92 7.83 ;
        RECT 0.02 7.57 0.28 7.83 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -7.75 0 1.25 0.6 ;
        RECT -0.45 0 -0.2 1.8 ;
        RECT -3.05 0 -2.65 1.8 ;
        RECT -6.3 0 -5.9 1.8 ;
      LAYER MET2 ;
        RECT -0.1 0.25 0.4 0.55 ;
        RECT -0.05 0.2 0.35 0.6 ;
        RECT -1.3 0.25 -0.8 0.55 ;
        RECT -1.25 0.2 -0.85 0.6 ;
        RECT -2.5 0.25 -2 0.55 ;
        RECT -2.45 0.2 -2.05 0.6 ;
        RECT -3.7 0.25 -3.2 0.55 ;
        RECT -3.65 0.2 -3.25 0.6 ;
        RECT -4.9 0.25 -4.4 0.55 ;
        RECT -4.85 0.2 -4.45 0.6 ;
        RECT -6.1 0.25 -5.6 0.55 ;
        RECT -6.05 0.2 -5.65 0.6 ;
        RECT -7.3 0.25 -6.8 0.55 ;
        RECT -7.25 0.2 -6.85 0.6 ;
      LAYER VIA12 ;
        RECT -7.18 0.27 -6.92 0.53 ;
        RECT -5.98 0.27 -5.72 0.53 ;
        RECT -4.78 0.27 -4.52 0.53 ;
        RECT -3.58 0.27 -3.32 0.53 ;
        RECT -2.38 0.27 -2.12 0.53 ;
        RECT -1.18 0.27 -0.92 0.53 ;
        RECT 0.02 0.27 0.28 0.53 ;
    END
  END VSS
  OBS
    LAYER MET2 ;
      RECT -1 3.45 -0.5 3.85 ;
      RECT -3.2 3.45 -2.8 3.85 ;
      RECT -7.4 3.45 -6.9 3.85 ;
      RECT -7.4 3.5 -0.5 3.8 ;
      RECT -1.25 4.75 -0.85 5.15 ;
      RECT -1.3 4.8 -0.8 5.1 ;
    LAYER VIA12 ;
      RECT -0.88 3.52 -0.62 3.78 ;
      RECT -1.18 4.82 -0.92 5.08 ;
      RECT -3.13 3.52 -2.87 3.78 ;
      RECT -7.28 3.52 -7.02 3.78 ;
    LAYER MET1 ;
      RECT -1.3 4.75 -1.05 7.15 ;
      RECT -1.3 4.75 -0.9 5.3 ;
      RECT -1.3 4.8 -0.8 5.1 ;
      RECT -1.3 4.8 0.05 5.05 ;
      RECT -0.25 2.05 0.05 5.05 ;
      RECT -1.3 2.05 0.05 2.3 ;
      RECT -1.3 0.95 -1.05 2.3 ;
      RECT -2.05 5.25 -1.8 7.15 ;
      RECT -1.8 1.95 -1.55 5.5 ;
      RECT -5.15 4.7 -4.65 5 ;
      RECT -5.05 2.55 -4.75 5 ;
      RECT -5.05 2.55 -1.55 2.85 ;
      RECT -2.05 0.95 -1.8 2.2 ;
      RECT -4.6 5.45 -4.35 7.15 ;
      RECT -6.6 5.45 -4.35 5.7 ;
      RECT -6.6 2.05 -6.35 5.7 ;
      RECT -6.65 4.15 -6.2 4.45 ;
      RECT -6.6 2.05 -4.35 2.3 ;
      RECT -4.6 0.95 -4.35 2.3 ;
      RECT -7.15 0.95 -6.9 7.15 ;
      RECT -7.25 3.45 -6.9 3.85 ;
      RECT -7.4 3.5 -6.9 3.8 ;
      RECT -7.3 3.45 -6.9 3.8 ;
      RECT -1 3.5 -0.5 3.8 ;
      RECT -3.25 3.5 -2.75 3.8 ;
  END
END gf180mcu_osu_sc_12T_dlatn_1
