* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

.option scale=0.05u

.subckt gf180mcu_osu_sc_gp9t3v3__tbuf_4 A Y EN EN_BAR
X0 Y a_17_19 VSS VSS nmos_3p3 w=17 l=6
X1 Y a_17_19 VSS VSS nmos_3p3 w=17 l=6
X2 Y a_17_19 VDD VDD pmos_3p3 w=34 l=6
X3 Y a_17_19 VDD VDD pmos_3p3 w=34 l=6
X4 a_33_19 EN a_17_19 VSS nmos_3p3 w=17 l=6
X5 VSS a_17_19 Y VSS nmos_3p3 w=17 l=6
X6 VSS a_17_19 Y VSS nmos_3p3 w=17 l=6
X7 a_33_70 EN_BAR a_17_19 VDD pmos_3p3 w=34 l=6
X8 VDD a_17_19 Y VDD pmos_3p3 w=34 l=6
X9 VSS A a_33_19 VSS nmos_3p3 w=17 l=6
X10 VDD a_17_19 Y VDD pmos_3p3 w=34 l=6
X11 VDD A a_33_70 VDD pmos_3p3 w=34 l=6
.ends

** hspice subcircuit dictionary
