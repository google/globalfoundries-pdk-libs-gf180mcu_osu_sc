# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_nand2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_nand2_1 0 -0.15 ;
  SIZE 3.1 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.6 3.35 1.1 3.65 ;
      LAYER MET2 ;
        RECT 0.6 3.3 1.1 3.7 ;
      LAYER VIA12 ;
        RECT 0.72 3.37 0.98 3.63 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 2.7 2.4 3 ;
      LAYER MET2 ;
        RECT 1.9 2.65 2.4 3.05 ;
      LAYER VIA12 ;
        RECT 2.02 2.72 2.28 2.98 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 3.1 7.95 ;
        RECT 2.25 5.3 2.5 7.95 ;
        RECT 0.55 5.3 0.8 7.95 ;
      LAYER MET2 ;
        RECT 1.65 7.4 2.15 7.7 ;
        RECT 1.7 7.35 2.1 7.75 ;
        RECT 0.45 7.4 0.95 7.7 ;
        RECT 0.5 7.35 0.9 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
        RECT 1.77 7.42 2.03 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 3.1 0.45 ;
        RECT 2.1 -0.15 2.35 1.65 ;
      LAYER MET2 ;
        RECT 1.65 0.1 2.15 0.4 ;
        RECT 1.7 0.05 2.1 0.45 ;
        RECT 0.45 0.1 0.95 0.4 ;
        RECT 0.5 0.05 0.9 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
        RECT 1.77 0.12 2.03 0.38 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.3 4 1.8 4.3 ;
        RECT 1.4 1.75 1.65 7 ;
        RECT 0.7 1.75 1.65 2 ;
        RECT 0.7 0.8 0.95 2 ;
      LAYER MET2 ;
        RECT 1.3 3.95 1.8 4.35 ;
      LAYER VIA12 ;
        RECT 1.42 4.02 1.68 4.28 ;
    END
  END Y
END gf180mcu_osu_sc_12T_nand2_1
