* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__addh_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__addh_1 A B S CO VDD VSS
X0 VDD B a_19_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_19_14# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD a_19_14# CO VDD pmos_3p3 w=1.7u l=0.3u
X3 a_19_14# B a_42_19# VSS nmos_3p3 w=0.85u l=0.3u
X4 S a_91_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X5 VSS a_19_14# CO VSS nmos_3p3 w=0.85u l=0.3u
X6 S a_91_19# VDD VDD pmos_3p3 w=1.7u l=0.3u
X7 a_91_19# B a_91_109# VDD pmos_3p3 w=1.7u l=0.3u
X8 VDD a_19_14# a_91_19# VDD pmos_3p3 w=1.7u l=0.3u
X9 a_91_109# A VDD VDD pmos_3p3 w=1.7u l=0.3u
X10 a_91_19# A a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X11 a_42_19# A VSS VSS nmos_3p3 w=0.85u l=0.3u
X12 VSS a_19_14# a_75_19# VSS nmos_3p3 w=0.85u l=0.3u
X13 a_75_19# B a_91_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
