# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai31_1 0 0 ;
  SIZE 4.9 BY 6.35 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 5.65 4.9 6.35 ;
        RECT 3.95 4.55 4.2 6.35 ;
        RECT 1 3.6 1.25 6.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.9 0.7 ;
        RECT 2.25 0 2.5 1.5 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 2.3 2.25 2.6 ;
      LAYER Metal2 ;
        RECT 1.75 2.25 2.25 2.65 ;
      LAYER Via1 ;
        RECT 1.87 2.32 2.13 2.58 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.55 2.95 3.05 3.25 ;
      LAYER Metal2 ;
        RECT 2.55 2.9 3.05 3.3 ;
      LAYER Via1 ;
        RECT 2.67 2.97 2.93 3.23 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.75 2.3 1.25 2.6 ;
      LAYER Metal2 ;
        RECT 0.75 2.25 1.25 2.65 ;
      LAYER Via1 ;
        RECT 0.87 2.32 1.13 2.58 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.25 2.3 3.75 2.6 ;
      LAYER Metal2 ;
        RECT 3.25 2.25 3.75 2.65 ;
      LAYER Via1 ;
        RECT 3.37 2.32 3.63 2.58 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 3.6 4.4 3.9 ;
        RECT 4 3.55 4.35 3.9 ;
        RECT 4.05 1.05 4.3 3.9 ;
        RECT 3 3.6 3.35 5.3 ;
      LAYER Metal2 ;
        RECT 3.9 3.6 4.4 3.9 ;
        RECT 3.95 3.55 4.35 3.95 ;
      LAYER Via1 ;
        RECT 4.02 3.62 4.28 3.88 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.75 3.45 2 ;
      RECT 3.1 1.05 3.45 2 ;
      RECT 1.4 1.05 1.65 2 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai31_1
