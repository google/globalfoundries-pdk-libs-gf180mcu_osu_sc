magic
tech gf180mcuC
timestamp 1659975453
<< nwell >>
rect -81 97 293 159
<< nmos >>
rect -62 16 -56 33
rect -27 16 -21 33
rect -10 16 -4 33
rect 1 16 7 33
rect 36 16 42 33
rect 52 16 58 33
rect 69 16 75 33
rect 80 16 86 33
rect 97 16 103 33
rect 108 16 114 33
rect 125 16 131 33
rect 136 16 142 33
rect 153 16 159 33
rect 188 16 194 33
rect 199 16 205 33
rect 216 16 222 33
rect 251 16 257 33
rect 268 16 274 33
<< pmos >>
rect -62 106 -56 140
rect -30 106 -24 140
rect -13 106 -7 140
rect 4 106 10 140
rect 36 106 42 140
rect 52 106 58 140
rect 69 106 75 140
rect 80 106 86 140
rect 97 106 103 140
rect 108 106 114 140
rect 125 106 131 140
rect 136 106 142 140
rect 153 106 159 140
rect 185 106 191 140
rect 202 106 208 140
rect 219 106 225 140
rect 251 106 257 140
rect 268 106 274 140
<< ndiff >>
rect -72 31 -62 33
rect -72 18 -70 31
rect -65 18 -62 31
rect -72 16 -62 18
rect -56 31 -46 33
rect -56 18 -53 31
rect -48 18 -46 31
rect -56 16 -46 18
rect -37 31 -27 33
rect -37 18 -35 31
rect -30 18 -27 31
rect -37 16 -27 18
rect -21 31 -10 33
rect -21 18 -18 31
rect -13 18 -10 31
rect -21 16 -10 18
rect -4 16 1 33
rect 7 31 17 33
rect 7 18 10 31
rect 15 18 17 31
rect 7 16 17 18
rect 26 31 36 33
rect 26 18 28 31
rect 33 18 36 31
rect 26 16 36 18
rect 42 16 52 33
rect 58 31 69 33
rect 58 18 61 31
rect 66 18 69 31
rect 58 16 69 18
rect 75 16 80 33
rect 86 23 97 33
rect 86 18 89 23
rect 94 18 97 23
rect 86 16 97 18
rect 103 16 108 33
rect 114 31 125 33
rect 114 18 117 31
rect 122 18 125 31
rect 114 16 125 18
rect 131 16 136 33
rect 142 31 153 33
rect 142 18 145 31
rect 150 18 153 31
rect 142 16 153 18
rect 159 31 169 33
rect 159 18 162 31
rect 167 18 169 31
rect 159 16 169 18
rect 178 31 188 33
rect 178 18 180 31
rect 185 18 188 31
rect 178 16 188 18
rect 194 16 199 33
rect 205 31 216 33
rect 205 18 208 31
rect 213 18 216 31
rect 205 16 216 18
rect 222 31 232 33
rect 222 18 225 31
rect 230 18 232 31
rect 222 16 232 18
rect 241 31 251 33
rect 241 18 243 31
rect 248 18 251 31
rect 241 16 251 18
rect 257 31 268 33
rect 257 18 260 31
rect 265 18 268 31
rect 257 16 268 18
rect 274 31 284 33
rect 274 18 277 31
rect 282 18 284 31
rect 274 16 284 18
<< pdiff >>
rect -72 138 -62 140
rect -72 108 -70 138
rect -65 108 -62 138
rect -72 106 -62 108
rect -56 138 -46 140
rect -56 108 -53 138
rect -48 108 -46 138
rect -56 106 -46 108
rect -40 138 -30 140
rect -40 108 -38 138
rect -33 108 -30 138
rect -40 106 -30 108
rect -24 138 -13 140
rect -24 123 -21 138
rect -16 123 -13 138
rect -24 106 -13 123
rect -7 138 4 140
rect -7 123 -4 138
rect 1 123 4 138
rect -7 106 4 123
rect 10 138 20 140
rect 10 123 13 138
rect 18 123 20 138
rect 10 106 20 123
rect 26 138 36 140
rect 26 108 28 138
rect 33 108 36 138
rect 26 106 36 108
rect 42 106 52 140
rect 58 138 69 140
rect 58 108 61 138
rect 66 108 69 138
rect 58 106 69 108
rect 75 106 80 140
rect 86 138 97 140
rect 86 108 89 138
rect 94 108 97 138
rect 86 106 97 108
rect 103 106 108 140
rect 114 138 125 140
rect 114 123 117 138
rect 122 123 125 138
rect 114 106 125 123
rect 131 106 136 140
rect 142 138 153 140
rect 142 123 145 138
rect 150 123 153 138
rect 142 106 153 123
rect 159 138 169 140
rect 159 108 162 138
rect 167 108 169 138
rect 159 106 169 108
rect 175 138 185 140
rect 175 124 177 138
rect 182 124 185 138
rect 175 106 185 124
rect 191 138 202 140
rect 191 133 194 138
rect 199 133 202 138
rect 191 106 202 133
rect 208 138 219 140
rect 208 125 211 138
rect 216 125 219 138
rect 208 106 219 125
rect 225 138 235 140
rect 225 108 228 138
rect 233 108 235 138
rect 225 106 235 108
rect 241 138 251 140
rect 241 108 243 138
rect 248 108 251 138
rect 241 106 251 108
rect 257 138 268 140
rect 257 108 260 138
rect 265 108 268 138
rect 257 106 268 108
rect 274 138 284 140
rect 274 108 277 138
rect 282 108 284 138
rect 274 106 284 108
<< ndiffc >>
rect -70 18 -65 31
rect -53 18 -48 31
rect -35 18 -30 31
rect -18 18 -13 31
rect 10 18 15 31
rect 28 18 33 31
rect 61 18 66 31
rect 89 18 94 23
rect 117 18 122 31
rect 145 18 150 31
rect 162 18 167 31
rect 180 18 185 31
rect 208 18 213 31
rect 225 18 230 31
rect 243 18 248 31
rect 260 18 265 31
rect 277 18 282 31
<< pdiffc >>
rect -70 108 -65 138
rect -53 108 -48 138
rect -38 108 -33 138
rect -21 123 -16 138
rect -4 123 1 138
rect 13 123 18 138
rect 28 108 33 138
rect 61 108 66 138
rect 89 108 94 138
rect 117 123 122 138
rect 145 123 150 138
rect 162 108 167 138
rect 177 124 182 138
rect 194 133 199 138
rect 211 125 216 138
rect 228 108 233 138
rect 243 108 248 138
rect 260 108 265 138
rect 277 108 282 138
<< psubdiff >>
rect -72 7 -63 9
rect -72 2 -70 7
rect -65 2 -63 7
rect -72 0 -63 2
rect -47 7 -38 9
rect -47 2 -45 7
rect -40 2 -38 7
rect -47 0 -38 2
rect -23 7 -14 9
rect -23 2 -21 7
rect -16 2 -14 7
rect -23 0 -14 2
rect 1 7 10 9
rect 1 2 3 7
rect 8 2 10 7
rect 1 0 10 2
rect 25 7 34 9
rect 25 2 27 7
rect 32 2 34 7
rect 25 0 34 2
rect 49 7 58 9
rect 49 2 51 7
rect 56 2 58 7
rect 49 0 58 2
rect 73 7 82 9
rect 73 2 75 7
rect 80 2 82 7
rect 73 0 82 2
rect 97 7 106 9
rect 97 2 99 7
rect 104 2 106 7
rect 97 0 106 2
rect 121 7 130 9
rect 121 2 123 7
rect 128 2 130 7
rect 121 0 130 2
rect 145 7 154 9
rect 145 2 147 7
rect 152 2 154 7
rect 145 0 154 2
rect 169 7 178 9
rect 169 2 171 7
rect 176 2 178 7
rect 169 0 178 2
rect 193 7 202 9
rect 193 2 195 7
rect 200 2 202 7
rect 193 0 202 2
rect 217 7 226 9
rect 217 2 219 7
rect 224 2 226 7
rect 217 0 226 2
rect 241 7 250 9
rect 241 2 243 7
rect 248 2 250 7
rect 241 0 250 2
rect 265 7 274 9
rect 265 2 267 7
rect 272 2 274 7
rect 265 0 274 2
<< nsubdiff >>
rect -72 154 -63 156
rect -72 149 -70 154
rect -65 149 -63 154
rect -72 147 -63 149
rect -47 154 -38 156
rect -47 149 -45 154
rect -40 149 -38 154
rect -47 147 -38 149
rect -23 154 -14 156
rect -23 149 -21 154
rect -16 149 -14 154
rect -23 147 -14 149
rect 1 154 10 156
rect 1 149 3 154
rect 8 149 10 154
rect 1 147 10 149
rect 25 154 34 156
rect 25 149 27 154
rect 32 149 34 154
rect 25 147 34 149
rect 49 154 58 156
rect 49 149 51 154
rect 56 149 58 154
rect 49 147 58 149
rect 73 154 82 156
rect 73 149 75 154
rect 80 149 82 154
rect 73 147 82 149
rect 97 154 106 156
rect 97 149 99 154
rect 104 149 106 154
rect 97 147 106 149
rect 121 154 130 156
rect 121 149 123 154
rect 128 149 130 154
rect 121 147 130 149
rect 145 154 154 156
rect 145 149 147 154
rect 152 149 154 154
rect 145 147 154 149
rect 169 154 178 156
rect 169 149 171 154
rect 176 149 178 154
rect 169 147 178 149
rect 193 154 202 156
rect 193 149 195 154
rect 200 149 202 154
rect 193 147 202 149
rect 217 154 226 156
rect 217 149 219 154
rect 224 149 226 154
rect 217 147 226 149
rect 241 154 250 156
rect 241 149 243 154
rect 248 149 250 154
rect 241 147 250 149
rect 265 154 274 156
rect 265 149 267 154
rect 272 149 274 154
rect 265 147 274 149
<< psubdiffcont >>
rect -70 2 -65 7
rect -45 2 -40 7
rect -21 2 -16 7
rect 3 2 8 7
rect 27 2 32 7
rect 51 2 56 7
rect 75 2 80 7
rect 99 2 104 7
rect 123 2 128 7
rect 147 2 152 7
rect 171 2 176 7
rect 195 2 200 7
rect 219 2 224 7
rect 243 2 248 7
rect 267 2 272 7
<< nsubdiffcont >>
rect -70 149 -65 154
rect -45 149 -40 154
rect -21 149 -16 154
rect 3 149 8 154
rect 27 149 32 154
rect 51 149 56 154
rect 75 149 80 154
rect 99 149 104 154
rect 123 149 128 154
rect 147 149 152 154
rect 171 149 176 154
rect 195 149 200 154
rect 219 149 224 154
rect 243 149 248 154
rect 267 149 272 154
<< polysilicon >>
rect -62 140 -56 145
rect -30 140 -24 145
rect -13 140 -7 145
rect 4 140 10 145
rect 36 140 42 145
rect 52 140 58 145
rect 69 140 75 145
rect 80 140 86 145
rect 97 140 103 145
rect 108 140 114 145
rect 125 140 131 145
rect 136 140 142 145
rect 153 140 159 145
rect 185 140 191 145
rect 202 140 208 145
rect 219 140 225 145
rect 251 140 257 145
rect 268 140 274 145
rect -62 101 -56 106
rect -69 99 -56 101
rect -69 94 -67 99
rect -62 94 -56 99
rect -69 92 -56 94
rect -62 33 -56 92
rect -30 75 -24 106
rect -13 88 -7 106
rect -13 86 -1 88
rect -13 80 -11 86
rect -5 80 -1 86
rect -13 78 -1 80
rect -30 73 -18 75
rect -30 67 -26 73
rect -20 67 -18 73
rect -30 65 -18 67
rect -30 60 -24 65
rect -30 56 -21 60
rect -27 33 -21 56
rect -13 42 -7 78
rect 4 75 10 106
rect 36 75 42 106
rect 52 88 58 106
rect 52 86 62 88
rect 52 80 54 86
rect 60 80 62 86
rect 52 78 62 80
rect 4 73 18 75
rect 4 67 9 73
rect 15 67 18 73
rect 4 65 18 67
rect 36 73 48 75
rect 36 67 40 73
rect 46 67 48 73
rect 36 65 48 67
rect 4 42 10 65
rect -13 38 -4 42
rect -10 33 -4 38
rect 1 38 10 42
rect 1 33 7 38
rect 36 33 42 65
rect 69 61 75 106
rect 80 101 86 106
rect 97 101 103 106
rect 80 99 103 101
rect 80 94 83 99
rect 81 93 83 94
rect 89 94 103 99
rect 89 93 91 94
rect 81 89 91 93
rect 108 61 114 106
rect 125 88 131 106
rect 121 86 131 88
rect 121 80 123 86
rect 129 80 131 86
rect 121 78 131 80
rect 136 75 142 106
rect 153 88 159 106
rect 153 86 163 88
rect 153 80 155 86
rect 161 80 163 86
rect 153 78 163 80
rect 135 73 145 75
rect 135 67 137 73
rect 143 67 145 73
rect 135 65 145 67
rect 121 61 131 62
rect 52 60 131 61
rect 52 55 123 60
rect 52 33 58 55
rect 121 54 123 55
rect 129 54 131 60
rect 121 52 131 54
rect 65 47 75 49
rect 81 47 91 49
rect 65 41 67 47
rect 73 41 75 47
rect 65 39 75 41
rect 69 33 75 39
rect 80 41 83 47
rect 89 41 103 47
rect 80 39 103 41
rect 80 33 86 39
rect 97 33 103 39
rect 108 46 118 48
rect 108 40 110 46
rect 116 40 118 46
rect 108 38 118 40
rect 108 33 114 38
rect 125 33 131 52
rect 136 33 142 65
rect 153 33 159 78
rect 185 48 191 106
rect 202 88 208 106
rect 196 86 208 88
rect 196 80 200 86
rect 206 80 208 86
rect 196 78 208 80
rect 177 46 191 48
rect 177 40 180 46
rect 186 42 191 46
rect 202 42 208 78
rect 219 60 225 106
rect 251 62 257 106
rect 268 88 274 106
rect 262 86 274 88
rect 262 80 264 86
rect 270 80 274 86
rect 262 78 274 80
rect 186 40 194 42
rect 177 38 194 40
rect 188 33 194 38
rect 199 38 208 42
rect 216 56 225 60
rect 245 60 257 62
rect 216 48 222 56
rect 245 54 249 60
rect 255 54 257 60
rect 245 52 257 54
rect 216 46 228 48
rect 216 40 220 46
rect 226 40 228 46
rect 216 38 228 40
rect 199 33 205 38
rect 216 33 222 38
rect 251 33 257 52
rect 268 33 274 78
rect -62 11 -56 16
rect -27 11 -21 16
rect -10 11 -4 16
rect 1 11 7 16
rect 36 11 42 16
rect 52 11 58 16
rect 69 11 75 16
rect 80 11 86 16
rect 97 11 103 16
rect 108 11 114 16
rect 125 11 131 16
rect 136 11 142 16
rect 153 11 159 16
rect 188 11 194 16
rect 199 11 205 16
rect 216 11 222 16
rect 251 11 257 16
rect 268 11 274 16
<< polycontact >>
rect -67 94 -62 99
rect -11 80 -5 86
rect -26 67 -20 73
rect 54 80 60 86
rect 9 67 15 73
rect 40 67 46 73
rect 83 93 89 99
rect 123 80 129 86
rect 155 80 161 86
rect 137 67 143 73
rect 123 54 129 60
rect 67 41 73 47
rect 83 41 89 47
rect 110 40 116 46
rect 200 80 206 86
rect 180 40 186 46
rect 264 80 270 86
rect 249 54 255 60
rect 220 40 226 46
<< metal1 >>
rect -81 154 293 159
rect -81 148 -70 154
rect -64 148 -46 154
rect -40 148 -22 154
rect -16 148 2 154
rect 8 148 26 154
rect 32 148 50 154
rect 56 148 74 154
rect 80 148 98 154
rect 104 148 122 154
rect 128 148 146 154
rect 152 148 170 154
rect 176 148 194 154
rect 200 148 218 154
rect 224 148 242 154
rect 248 148 266 154
rect 272 148 293 154
rect -81 147 293 148
rect -70 138 -65 147
rect -70 106 -65 108
rect -53 138 -48 140
rect -70 93 -68 99
rect -62 93 -60 99
rect -53 47 -48 108
rect -38 138 -33 140
rect -21 138 -16 140
rect -21 116 -16 123
rect -4 138 1 147
rect -4 121 1 123
rect 13 138 18 140
rect 13 116 18 123
rect -21 111 18 116
rect 28 138 33 147
rect -38 52 -33 108
rect 28 106 33 108
rect 61 138 66 140
rect 61 101 66 108
rect 89 138 94 147
rect 117 138 122 140
rect 117 121 122 123
rect 145 138 150 147
rect 145 121 150 123
rect 162 138 167 140
rect 89 106 94 108
rect 99 116 122 121
rect 28 96 66 101
rect -13 80 -11 86
rect -5 80 -3 86
rect 28 73 33 96
rect 81 93 83 99
rect 89 93 91 99
rect 52 80 54 86
rect 60 80 67 86
rect 73 80 75 86
rect -28 67 -26 73
rect -20 67 -18 73
rect 7 67 9 73
rect 15 67 33 73
rect 38 67 40 73
rect 46 67 48 73
rect -38 47 -13 52
rect 9 47 14 48
rect 28 47 33 67
rect 67 47 73 80
rect 83 47 89 93
rect 99 71 104 116
rect 177 138 182 140
rect 194 138 199 147
rect 194 131 199 133
rect 211 138 216 140
rect 182 125 211 126
rect 182 124 216 125
rect 177 121 216 124
rect 228 138 233 140
rect 134 93 136 99
rect 142 93 144 99
rect 162 97 167 108
rect 180 99 186 101
rect 228 99 233 108
rect 243 138 248 140
rect 98 66 104 71
rect 110 80 123 86
rect 129 80 131 86
rect -55 41 -53 47
rect -47 41 -45 47
rect -18 41 9 47
rect 15 41 17 47
rect 28 42 48 47
rect -53 40 -47 41
rect -70 31 -65 33
rect -70 9 -65 18
rect -53 31 -48 40
rect -53 16 -48 18
rect -35 31 -30 33
rect -35 9 -30 18
rect -18 31 -13 41
rect 9 40 14 41
rect 40 33 48 42
rect 65 41 67 47
rect 73 41 75 47
rect 81 41 83 47
rect 89 41 91 47
rect 98 34 103 66
rect 110 46 116 80
rect 136 73 142 93
rect 162 92 173 97
rect 153 80 155 86
rect 161 80 163 86
rect 168 73 173 92
rect 186 93 228 99
rect 234 93 236 99
rect 180 91 186 93
rect 198 80 200 86
rect 206 80 208 86
rect 135 67 137 73
rect 143 67 145 73
rect 162 68 173 73
rect 162 60 168 68
rect 228 60 233 93
rect 243 86 248 108
rect 260 138 265 147
rect 260 106 265 108
rect 277 138 282 140
rect 277 100 282 108
rect 277 99 287 100
rect 277 93 279 99
rect 285 93 287 99
rect 277 92 286 93
rect 243 80 264 86
rect 270 80 272 86
rect 121 54 123 60
rect 129 54 131 60
rect 162 52 168 54
rect 208 54 249 60
rect 255 54 257 60
rect 108 40 110 46
rect 116 40 118 46
rect -18 16 -13 18
rect 10 31 15 33
rect 10 9 15 18
rect 28 31 33 33
rect 40 31 66 33
rect 40 28 61 31
rect 28 9 33 18
rect 98 29 117 34
rect 123 28 125 34
rect 145 31 150 33
rect 61 16 66 18
rect 89 23 94 25
rect 89 9 94 18
rect 117 16 122 18
rect 145 9 150 18
rect 162 31 167 52
rect 178 40 180 46
rect 186 40 188 46
rect 162 16 167 18
rect 180 31 185 33
rect 180 9 185 18
rect 208 31 213 54
rect 218 40 220 46
rect 226 40 228 46
rect 265 43 270 80
rect 243 38 270 43
rect 208 16 213 18
rect 225 31 230 33
rect 225 9 230 18
rect 243 31 248 38
rect 243 16 248 18
rect 260 31 265 33
rect 260 9 265 18
rect 277 31 282 92
rect 277 16 282 18
rect -81 8 293 9
rect -81 2 -70 8
rect -64 2 -46 8
rect -40 2 -22 8
rect -16 2 2 8
rect 8 2 26 8
rect 32 2 50 8
rect 56 2 74 8
rect 80 2 98 8
rect 104 2 122 8
rect 128 2 146 8
rect 152 2 170 8
rect 176 2 194 8
rect 200 2 218 8
rect 224 2 242 8
rect 248 2 266 8
rect 272 2 293 8
rect -81 -3 293 2
<< via1 >>
rect -70 149 -65 154
rect -65 149 -64 154
rect -70 148 -64 149
rect -46 149 -45 154
rect -45 149 -40 154
rect -46 148 -40 149
rect -22 149 -21 154
rect -21 149 -16 154
rect -22 148 -16 149
rect 2 149 3 154
rect 3 149 8 154
rect 2 148 8 149
rect 26 149 27 154
rect 27 149 32 154
rect 26 148 32 149
rect 50 149 51 154
rect 51 149 56 154
rect 50 148 56 149
rect 74 149 75 154
rect 75 149 80 154
rect 74 148 80 149
rect 98 149 99 154
rect 99 149 104 154
rect 98 148 104 149
rect 122 149 123 154
rect 123 149 128 154
rect 122 148 128 149
rect 146 149 147 154
rect 147 149 152 154
rect 146 148 152 149
rect 170 149 171 154
rect 171 149 176 154
rect 170 148 176 149
rect 194 149 195 154
rect 195 149 200 154
rect 194 148 200 149
rect 218 149 219 154
rect 219 149 224 154
rect 218 148 224 149
rect 242 149 243 154
rect 243 149 248 154
rect 242 148 248 149
rect 266 149 267 154
rect 267 149 272 154
rect 266 148 272 149
rect -68 94 -67 99
rect -67 94 -62 99
rect -68 93 -62 94
rect -11 80 -5 86
rect 67 80 73 86
rect -26 67 -20 73
rect 9 67 15 73
rect 40 67 46 73
rect 136 93 142 99
rect 123 80 129 86
rect -53 41 -47 47
rect 9 41 15 47
rect 83 41 89 47
rect 155 80 161 86
rect 180 93 186 99
rect 228 93 234 99
rect 200 80 206 86
rect 137 67 143 73
rect 279 93 285 99
rect 264 80 270 86
rect 123 54 129 60
rect 162 54 168 60
rect 249 54 255 60
rect 117 31 123 34
rect 117 28 122 31
rect 122 28 123 31
rect 180 40 186 46
rect 220 40 226 46
rect -70 7 -64 8
rect -70 2 -65 7
rect -65 2 -64 7
rect -46 7 -40 8
rect -46 2 -45 7
rect -45 2 -40 7
rect -22 7 -16 8
rect -22 2 -21 7
rect -21 2 -16 7
rect 2 7 8 8
rect 2 2 3 7
rect 3 2 8 7
rect 26 7 32 8
rect 26 2 27 7
rect 27 2 32 7
rect 50 7 56 8
rect 50 2 51 7
rect 51 2 56 7
rect 74 7 80 8
rect 74 2 75 7
rect 75 2 80 7
rect 98 7 104 8
rect 98 2 99 7
rect 99 2 104 7
rect 122 7 128 8
rect 122 2 123 7
rect 123 2 128 7
rect 146 7 152 8
rect 146 2 147 7
rect 147 2 152 7
rect 170 7 176 8
rect 170 2 171 7
rect 171 2 176 7
rect 194 7 200 8
rect 194 2 195 7
rect 195 2 200 7
rect 218 7 224 8
rect 218 2 219 7
rect 219 2 224 7
rect 242 7 248 8
rect 242 2 243 7
rect 243 2 248 7
rect 266 7 272 8
rect 266 2 267 7
rect 267 2 272 7
<< metal2 >>
rect -71 154 -63 155
rect -47 154 -39 155
rect -23 154 -15 155
rect 1 154 9 155
rect 25 154 33 155
rect 49 154 57 155
rect 73 154 81 155
rect 97 154 105 155
rect 121 154 129 155
rect 145 154 153 155
rect 169 154 177 155
rect 193 154 201 155
rect 217 154 225 155
rect 241 154 249 155
rect 265 154 273 155
rect -72 148 -70 154
rect -64 148 -62 154
rect -48 148 -46 154
rect -40 148 -38 154
rect -24 148 -22 154
rect -16 148 -14 154
rect 0 148 2 154
rect 8 148 10 154
rect 24 148 26 154
rect 32 148 34 154
rect 48 148 50 154
rect 56 148 58 154
rect 72 148 74 154
rect 80 148 82 154
rect 96 148 98 154
rect 104 148 106 154
rect 120 148 122 154
rect 128 148 130 154
rect 144 148 146 154
rect 152 148 154 154
rect 168 148 170 154
rect 176 148 178 154
rect 192 148 194 154
rect 200 148 202 154
rect 216 148 218 154
rect 224 148 226 154
rect 240 148 242 154
rect 248 148 250 154
rect 264 148 266 154
rect 272 148 274 154
rect -71 147 -63 148
rect -47 147 -39 148
rect -23 147 -15 148
rect 1 147 9 148
rect 25 147 33 148
rect 49 147 57 148
rect 73 147 81 148
rect 97 147 105 148
rect 121 147 129 148
rect 145 147 153 148
rect 169 147 177 148
rect 193 147 201 148
rect 217 147 225 148
rect 241 147 249 148
rect 265 147 273 148
rect -11 106 206 112
rect -70 99 -60 100
rect -70 93 -68 99
rect -62 93 -60 99
rect -70 92 -60 93
rect -11 87 -5 106
rect 135 99 143 100
rect 179 99 187 100
rect 134 93 136 99
rect 142 93 180 99
rect 186 93 188 99
rect 135 92 143 93
rect 179 92 187 93
rect 200 87 206 106
rect 226 99 236 100
rect 278 99 286 100
rect 226 93 228 99
rect 234 93 236 99
rect 277 93 279 99
rect 285 93 287 99
rect 226 92 236 93
rect 278 92 286 93
rect -13 86 -3 87
rect -13 80 -11 86
rect -5 80 -3 86
rect -13 79 -3 80
rect 65 86 74 87
rect 121 86 131 87
rect 154 86 162 87
rect 198 86 208 87
rect 263 86 271 87
rect 65 80 67 86
rect 73 80 123 86
rect 129 80 155 86
rect 161 80 163 86
rect 198 80 200 86
rect 206 80 208 86
rect 262 80 264 86
rect 270 80 272 86
rect 65 79 74 80
rect 121 79 131 80
rect 154 79 162 80
rect 198 79 208 80
rect 263 79 271 80
rect -28 73 -18 74
rect -28 67 -26 73
rect -20 67 -18 73
rect -28 66 -18 67
rect 7 73 17 74
rect 7 67 9 73
rect 15 67 17 73
rect 7 66 17 67
rect 38 73 48 74
rect 136 73 144 74
rect 38 67 40 73
rect 46 67 48 73
rect 135 67 137 73
rect 143 67 145 73
rect 38 66 48 67
rect 136 66 144 67
rect -55 47 -45 48
rect -26 47 -20 66
rect 122 60 130 61
rect 161 60 169 61
rect 248 60 256 61
rect 121 54 123 60
rect 129 54 162 60
rect 168 54 171 60
rect 241 54 249 60
rect 255 54 257 60
rect 122 53 130 54
rect 161 53 169 54
rect 248 53 256 54
rect -55 41 -53 47
rect -47 41 -20 47
rect -55 40 -45 41
rect -26 21 -20 41
rect 7 47 17 48
rect 82 47 90 48
rect 7 41 9 47
rect 15 41 83 47
rect 89 41 91 47
rect 178 46 188 47
rect 7 40 17 41
rect 82 40 90 41
rect 178 40 180 46
rect 186 40 188 46
rect 178 39 188 40
rect 216 46 228 47
rect 216 40 220 46
rect 226 40 228 46
rect 216 39 228 40
rect 116 34 124 35
rect 178 34 186 39
rect 115 28 117 34
rect 123 28 186 34
rect 116 27 124 28
rect 216 21 222 39
rect -26 15 222 21
rect -71 8 -63 9
rect -47 8 -39 9
rect -23 8 -15 9
rect 1 8 9 9
rect 25 8 33 9
rect 49 8 57 9
rect 73 8 81 9
rect 97 8 105 9
rect 121 8 129 9
rect 145 8 153 9
rect 169 8 177 9
rect 193 8 201 9
rect 217 8 225 9
rect 241 8 249 9
rect 265 8 273 9
rect -72 2 -70 8
rect -64 2 -62 8
rect -48 2 -46 8
rect -40 2 -38 8
rect -24 2 -22 8
rect -16 2 -14 8
rect 0 2 2 8
rect 8 2 10 8
rect 24 2 26 8
rect 32 2 34 8
rect 48 2 50 8
rect 56 2 58 8
rect 72 2 74 8
rect 80 2 82 8
rect 96 2 98 8
rect 104 2 106 8
rect 120 2 122 8
rect 128 2 130 8
rect 144 2 146 8
rect 152 2 154 8
rect 168 2 170 8
rect 176 2 178 8
rect 192 2 194 8
rect 200 2 202 8
rect 216 2 218 8
rect 224 2 226 8
rect 240 2 242 8
rect 248 2 250 8
rect 264 2 266 8
rect 272 2 274 8
rect -71 1 -63 2
rect -47 1 -39 2
rect -23 1 -15 2
rect 1 1 9 2
rect 25 1 33 2
rect 49 1 57 2
rect 73 1 81 2
rect 97 1 105 2
rect 121 1 129 2
rect 145 1 153 2
rect 169 1 177 2
rect 193 1 201 2
rect 217 1 225 2
rect 241 1 249 2
rect 265 1 273 2
<< labels >>
rlabel metal2 43 70 43 70 1 D
port 1 n
rlabel metal2 282 96 282 96 1 Q
port 5 n
rlabel metal2 -67 151 -67 151 1 VDD
rlabel metal2 -67 4 -67 4 1 GND
rlabel metal2 -65 96 -65 96 1 RN
port 4 n
rlabel metal2 203 83 203 83 1 SN
port 3 n
rlabel metal2 267 83 267 83 1 QN
port 8 n
rlabel metal2 158 83 158 83 1 CLK
port 9 n
<< end >>
