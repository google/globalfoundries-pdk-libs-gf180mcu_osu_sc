magic
tech gf180mcuC
timestamp 1659966734
<< nwell >>
rect 0 97 176 159
<< metal1 >>
rect 0 147 176 159
rect 0 -3 176 9
<< labels >>
rlabel metal1 8 153 8 153 1 VDD
rlabel metal1 7 2 7 2 1 GND
<< end >>
