# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__aoi31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__aoi31_1 0 0 ;
  SIZE 4.95 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.95 6.15 ;
        RECT 2.25 4.25 2.5 6.15 ;
        RECT 0.55 3.75 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.95 0.6 ;
        RECT 3.8 0 4.05 1.8 ;
        RECT 0.95 0 1.2 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.6 2.85 2.1 3.15 ;
      LAYER MET2 ;
        RECT 1.6 2.8 2.1 3.2 ;
      LAYER VIA12 ;
        RECT 1.72 2.87 1.98 3.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.5 2.85 3 3.15 ;
      LAYER MET2 ;
        RECT 2.5 2.8 3 3.2 ;
      LAYER VIA12 ;
        RECT 2.62 2.87 2.88 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 2.85 1.25 3.15 ;
      LAYER MET2 ;
        RECT 0.75 2.8 1.25 3.2 ;
      LAYER VIA12 ;
        RECT 0.87 2.87 1.13 3.13 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.35 2.75 3.65 3.25 ;
      LAYER MET2 ;
        RECT 3.3 2.75 3.7 3.25 ;
      LAYER VIA12 ;
        RECT 3.37 2.87 3.63 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.95 2.25 4.45 2.5 ;
        RECT 3.95 2.2 4.45 2.5 ;
        RECT 4.05 2.15 4.3 2.55 ;
        RECT 3.95 2.2 4.2 5.2 ;
        RECT 2.95 0.95 3.2 2.5 ;
      LAYER MET2 ;
        RECT 4 2.1 4.4 2.6 ;
      LAYER VIA12 ;
        RECT 4.07 2.22 4.33 2.48 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 3.1 3.75 3.35 5.2 ;
      RECT 1.4 3.75 1.65 5.2 ;
      RECT 1.4 3.75 3.35 4 ;
  END
END gf180mcu_osu_sc_gp9t3v3__aoi31_1
