magic
tech gf180mcuC
timestamp 1661875002
<< error_p >>
rect 0 111 18 123
rect 4 61 18 111
rect 0 0 5 12
<< nwell >>
rect 0 61 4 123
<< metal1 >>
rect 0 111 4 123
rect 0 0 4 12
<< labels >>
rlabel metal1 2 116 2 116 3 VDD
rlabel metal1 2 5 2 5 2 GND
<< end >>
