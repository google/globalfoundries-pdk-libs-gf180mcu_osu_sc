# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__oai21_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai21_1 0 0 ;
  SIZE 3.9 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.9 8.1 ;
        RECT 2.95 5.45 3.2 8.1 ;
        RECT 0.65 5.45 0.9 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.9 0.6 ;
        RECT 1.35 0 1.6 1.5 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.45 3.5 0.95 3.8 ;
      LAYER MET2 ;
        RECT 0.45 3.45 0.95 3.85 ;
      LAYER VIA12 ;
        RECT 0.57 3.52 0.83 3.78 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4.15 1.95 4.45 ;
      LAYER MET2 ;
        RECT 1.45 4.1 1.95 4.5 ;
      LAYER VIA12 ;
        RECT 1.57 4.17 1.83 4.43 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.2 3.5 2.7 3.8 ;
      LAYER MET2 ;
        RECT 2.2 3.45 2.7 3.85 ;
      LAYER VIA12 ;
        RECT 2.32 3.52 2.58 3.78 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.1 4.8 3.35 5.1 ;
        RECT 3.05 0.95 3.3 2.5 ;
        RECT 2.95 2.25 3.2 5.1 ;
        RECT 2.1 4.8 2.35 7.15 ;
      LAYER MET2 ;
        RECT 2.85 4.75 3.35 5.15 ;
      LAYER VIA12 ;
        RECT 2.97 4.82 3.23 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.5 1.75 2.45 2 ;
      RECT 2.2 0.95 2.45 2 ;
      RECT 0.5 0.95 0.75 2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai21_1
