* NGSPICE file created from gf180mcu_osu_sc_12T_aoi21_1.ext - technology: gf180mcuC

.inc "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/design.hspice"
.lib "/import/yukari1/lrburle/globalfoundries-pdk-libs-gf180mcu_osu_sc/char/techfiles/sm141064.hspice" typical

X0 Y B a_9_106# VDD pmos_3p3 w=1.7u l=0.3u
X1 a_9_106# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X2 VDD A0 a_9_106# VDD pmos_3p3 w=1.7u l=0.3u
X3 GND B Y GND nmos_3p3 w=0.85u l=0.3u
X4 a_28_16# A0 GND GND nmos_3p3 w=0.85u l=0.3u
X5 Y A1 a_28_16# GND nmos_3p3 w=0.85u l=0.3u
