# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_clkbuf_16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_clkbuf_16 0 0 ;
  SIZE 15.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 15.8 8.1 ;
        RECT 15 5.45 15.25 8.1 ;
        RECT 13.3 5.45 13.55 8.1 ;
        RECT 11.6 5.45 11.85 8.1 ;
        RECT 9.9 5.45 10.15 8.1 ;
        RECT 8.2 5.45 8.45 8.1 ;
        RECT 6.5 5.45 6.75 8.1 ;
        RECT 4.8 5.45 5.05 8.1 ;
        RECT 3.1 5.45 3.35 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 15.8 0.6 ;
        RECT 15 0 15.25 1.8 ;
        RECT 13.3 0 13.55 1.8 ;
        RECT 11.6 0 11.85 1.8 ;
        RECT 9.9 0 10.15 1.8 ;
        RECT 8.2 0 8.45 1.8 ;
        RECT 6.5 0 6.75 1.8 ;
        RECT 4.8 0 5.05 1.8 ;
        RECT 3.1 0 3.35 1.8 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 4.15 1.55 4.45 ;
      LAYER MET2 ;
        RECT 1.05 4.15 1.55 4.45 ;
        RECT 1.1 4.1 1.5 4.5 ;
      LAYER VIA12 ;
        RECT 1.17 4.17 1.43 4.43 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 4.85 14.55 5.15 ;
        RECT 14.15 0.95 14.4 7.15 ;
        RECT 2.25 2.05 14.4 2.3 ;
        RECT 12.45 0.95 12.7 7.15 ;
        RECT 10.75 0.95 11 7.15 ;
        RECT 9.05 0.95 9.3 7.15 ;
        RECT 7.35 0.95 7.6 7.15 ;
        RECT 5.65 0.95 5.9 7.15 ;
        RECT 3.95 0.95 4.2 7.15 ;
        RECT 2.25 0.95 2.5 7.15 ;
      LAYER MET2 ;
        RECT 14.05 4.8 14.55 5.2 ;
        RECT 14 4.85 14.55 5.15 ;
      LAYER VIA12 ;
        RECT 14.17 4.87 14.43 5.13 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 7.15 ;
      RECT 0.55 2.9 2 3.2 ;
  END
END gf180mcu_osu_sc_12T_clkbuf_16
