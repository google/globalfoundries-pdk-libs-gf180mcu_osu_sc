magic
tech gf180mcuC
timestamp 1661874473
<< nwell >>
rect 0 61 78 123
<< nmos >>
rect 22 19 28 36
rect 33 19 39 36
rect 50 19 56 36
<< pmos >>
rect 19 70 25 104
rect 36 70 42 104
rect 53 70 59 104
<< ndiff >>
rect 12 34 22 36
rect 12 21 14 34
rect 19 21 22 34
rect 12 19 22 21
rect 28 19 33 36
rect 39 31 50 36
rect 39 21 42 31
rect 47 21 50 31
rect 39 19 50 21
rect 56 26 66 36
rect 56 21 59 26
rect 64 21 66 26
rect 56 19 66 21
<< pdiff >>
rect 9 102 19 104
rect 9 87 11 102
rect 16 87 19 102
rect 9 70 19 87
rect 25 102 36 104
rect 25 87 28 102
rect 33 87 36 102
rect 25 70 36 87
rect 42 102 53 104
rect 42 87 45 102
rect 50 87 53 102
rect 42 70 53 87
rect 59 102 69 104
rect 59 88 62 102
rect 67 88 69 102
rect 59 70 69 88
<< ndiffc >>
rect 14 21 19 34
rect 42 21 47 31
rect 59 21 64 26
<< pdiffc >>
rect 11 87 16 102
rect 28 87 33 102
rect 45 87 50 102
rect 62 88 67 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
<< polysilicon >>
rect 19 104 25 109
rect 36 104 42 109
rect 53 104 59 109
rect 19 52 25 70
rect 36 65 42 70
rect 30 63 42 65
rect 30 57 34 63
rect 40 57 42 63
rect 30 55 42 57
rect 11 50 25 52
rect 11 44 14 50
rect 20 44 25 50
rect 11 43 25 44
rect 36 43 42 55
rect 53 52 59 70
rect 11 42 28 43
rect 19 39 28 42
rect 22 36 28 39
rect 33 38 42 43
rect 47 50 59 52
rect 47 44 49 50
rect 55 44 59 50
rect 47 42 59 44
rect 33 36 39 38
rect 50 36 56 42
rect 22 14 28 19
rect 33 14 39 19
rect 50 14 56 19
<< polycontact >>
rect 34 57 40 63
rect 14 44 20 50
rect 49 44 55 50
<< metal1 >>
rect 0 118 78 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 78 118
rect 0 111 78 112
rect 11 102 16 104
rect 11 80 16 87
rect 28 102 33 111
rect 28 85 33 87
rect 45 102 50 104
rect 45 80 50 87
rect 11 75 50 80
rect 62 102 67 104
rect 62 76 67 88
rect 60 70 62 76
rect 68 70 70 76
rect 32 57 34 63
rect 40 57 42 63
rect 12 44 14 50
rect 20 44 22 50
rect 47 44 49 50
rect 55 44 57 50
rect 62 38 67 70
rect 14 34 19 36
rect 14 12 19 21
rect 42 33 67 38
rect 42 31 47 33
rect 42 19 47 21
rect 59 26 64 28
rect 59 12 64 21
rect 0 11 78 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 78 11
rect 0 0 78 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 62 70 68 76
rect 34 57 40 63
rect 14 44 20 50
rect 49 44 55 50
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 11 118
rect 17 112 19 118
rect 33 112 35 118
rect 41 112 43 118
rect 57 112 59 118
rect 65 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 60 76 70 77
rect 60 70 62 76
rect 68 70 70 76
rect 60 69 70 70
rect 32 63 42 64
rect 32 57 34 63
rect 40 57 42 63
rect 32 56 42 57
rect 12 50 22 51
rect 12 44 14 50
rect 20 44 22 50
rect 12 43 22 44
rect 47 50 57 51
rect 47 44 49 50
rect 55 44 57 50
rect 47 43 57 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 11 11
rect 17 5 19 11
rect 33 5 35 11
rect 41 5 43 11
rect 57 5 59 11
rect 65 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 14 115 14 115 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 17 47 17 47 1 A0
port 5 n
rlabel metal2 37 60 37 60 1 A1
port 6 n
rlabel metal2 52 47 52 47 1 B
port 7 n
rlabel metal2 65 73 65 73 1 Y
port 4 n
<< end >>
