VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_9T_buf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_9T_buf_1 0 0 ;
  SIZE 3.2 BY 6.15 ;
  SYMMETRY X Y ;
  SITE 9T ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.05 2.85 1.55 3.15 ;
      LAYER MET2 ;
        RECT 1.05 2.85 1.55 3.15 ;
        RECT 1.1 2.8 1.5 3.2 ;
      LAYER VIA12 ;
        RECT 1.17 2.87 1.43 3.13 ;
    END
  END A
  PIN GND
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.2 0.6 ;
        RECT 1.4 0 1.75 1.8 ;
      LAYER MET2 ;
        RECT 1.65 0.25 2.15 0.55 ;
        RECT 1.7 0.2 2.1 0.6 ;
        RECT 0.45 0.25 0.95 0.55 ;
        RECT 0.5 0.2 0.9 0.6 ;
      LAYER VIA12 ;
        RECT 0.57 0.27 0.83 0.53 ;
        RECT 1.77 0.27 2.03 0.53 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 3.2 6.15 ;
        RECT 1.4 3.5 1.75 6.15 ;
      LAYER MET2 ;
        RECT 1.65 5.6 2.15 5.9 ;
        RECT 1.7 5.55 2.1 5.95 ;
        RECT 0.45 5.6 0.95 5.9 ;
        RECT 0.5 5.55 0.9 5.95 ;
      LAYER VIA12 ;
        RECT 0.57 5.62 0.83 5.88 ;
        RECT 1.77 5.62 2.03 5.88 ;
    END
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.25 1.5 2.75 1.8 ;
        RECT 2.35 0.95 2.6 1.8 ;
        RECT 2.25 3.5 2.75 3.8 ;
        RECT 2.35 3.5 2.6 5.2 ;
      LAYER MET2 ;
        RECT 2.25 3.45 2.75 3.85 ;
        RECT 2.25 1.45 2.75 1.85 ;
        RECT 2.35 1.45 2.65 3.85 ;
      LAYER VIA12 ;
        RECT 2.37 3.52 2.63 3.78 ;
        RECT 2.37 1.52 2.63 1.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 0.55 0.95 0.8 5.2 ;
      RECT 0.55 2.15 2.2 2.45 ;
  END
END gf180mcu_osu_sc_9T_buf_1
