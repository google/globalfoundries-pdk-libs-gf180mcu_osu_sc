# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__mux2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__mux2_1 0 0 ;
  SIZE 4.8 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 4.8 8.3 ;
        RECT 0.55 5.55 0.8 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 4.8 0.7 ;
        RECT 0.55 0 0.8 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.25 3.55 2.85 3.95 ;
        RECT 2.25 1.05 2.5 7.25 ;
      LAYER Metal2 ;
        RECT 2.35 3.55 2.85 3.95 ;
      LAYER Via1 ;
        RECT 2.47 3.62 2.73 3.88 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.75 4.2 4.25 4.6 ;
        RECT 3.95 1.05 4.2 7.25 ;
      LAYER Metal2 ;
        RECT 3.75 4.2 4.25 4.6 ;
      LAYER Via1 ;
        RECT 3.87 4.27 4.13 4.53 ;
    END
  END B
  PIN Sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.55 2.95 1.05 3.25 ;
      LAYER Metal2 ;
        RECT 0.55 2.9 1.05 3.3 ;
      LAYER Via1 ;
        RECT 0.67 2.97 0.93 3.23 ;
    END
  END Sel
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 4.85 3.5 5.25 ;
        RECT 3.1 1.05 3.35 7.25 ;
      LAYER Metal2 ;
        RECT 3 4.85 3.5 5.25 ;
      LAYER Via1 ;
        RECT 3.12 4.92 3.38 5.18 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      RECT 1.4 1.05 1.65 7.25 ;
      RECT 1.4 4.25 2 4.55 ;
      RECT 1.4 2.3 2 2.6 ;
  END
END gf180mcu_osu_sc_gp12t3v3__mux2_1
