# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__tinv_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tinv_1 0 0 ;
  SIZE 3.65 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 3.65 8.1 ;
        RECT 1.4 5.45 1.65 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 3.65 0.6 ;
        RECT 1.4 0 1.65 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.45 4.8 1.95 5.1 ;
      LAYER MET2 ;
        RECT 1.45 4.75 1.95 5.15 ;
      LAYER VIA12 ;
        RECT 1.57 4.82 1.83 5.08 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.7 2.2 3.2 2.5 ;
        RECT 1 2.2 1.5 2.5 ;
      LAYER MET2 ;
        RECT 2.7 2.15 3.2 2.55 ;
        RECT 1 2.2 3.2 2.5 ;
        RECT 1 2.15 1.5 2.55 ;
      LAYER VIA12 ;
        RECT 1.12 2.22 1.38 2.48 ;
        RECT 2.82 2.22 3.08 2.48 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 5.45 3.05 7.15 ;
        RECT 2.2 1.55 3.05 1.8 ;
        RECT 2.8 0.95 3.05 1.8 ;
        RECT 2.2 5.45 3.05 5.7 ;
        RECT 2.05 3.5 2.6 3.8 ;
        RECT 2.2 1.55 2.45 5.7 ;
      LAYER MET2 ;
        RECT 2.05 3.45 2.55 3.85 ;
      LAYER VIA12 ;
        RECT 2.17 3.52 2.43 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 2.7 4.75 3.2 5.15 ;
      RECT 2.8 4.15 3.1 5.15 ;
      RECT 0.35 4.1 0.85 4.5 ;
      RECT 0.35 4.15 3.1 4.45 ;
    LAYER VIA12 ;
      RECT 2.82 4.82 3.08 5.08 ;
      RECT 0.47 4.17 0.73 4.43 ;
    LAYER MET1 ;
      RECT 0.55 5.45 0.8 7.15 ;
      RECT 0.5 1.8 0.75 5.7 ;
      RECT 0.35 4.15 0.85 4.45 ;
      RECT 0.55 0.95 0.8 2.05 ;
      RECT 2.7 4.8 3.2 5.1 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tinv_1
