* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffr_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffr_1 D Q QN CLK RN VDD VSS
X0 a_122_16# CLK VDD VDD pfet_03p3 w=1.7u l=0.3u
X1 VDD a_205_70# a_201_111# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_62_100# CLK a_112_111# VDD pfet_03p3 w=1.7u l=0.3u
X3 a_145_111# a_122_16# a_62_100# VDD pfet_03p3 w=1.7u l=0.3u
X4 a_145_21# CLK a_62_100# VSS nfet_03p3 w=0.85u l=0.3u
X5 a_25_21# RN VDD VDD pfet_03p3 w=1.7u l=0.3u
X6 a_41_111# a_25_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X7 a_62_100# a_122_16# a_112_21# VSS nfet_03p3 w=0.85u l=0.3u
X8 a_112_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X9 a_205_70# a_184_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_25_21# RN VSS VSS nfet_03p3 w=0.85u l=0.3u
X11 VDD a_205_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X12 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X13 a_201_21# a_122_16# a_184_21# VSS nfet_03p3 w=0.85u l=0.3u
X14 VSS a_205_70# a_201_21# VSS nfet_03p3 w=0.85u l=0.3u
X15 a_205_70# a_25_21# a_273_111# VDD pfet_03p3 w=1.7u l=0.3u
X16 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X17 VSS a_205_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X18 a_273_111# a_184_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X19 VDD a_62_100# a_57_111# VDD pfet_03p3 w=1.7u l=0.3u
X20 VSS a_62_100# a_41_111# VSS nfet_03p3 w=0.85u l=0.3u
X21 a_112_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 a_57_111# a_25_21# a_41_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_173_21# a_41_111# VSS VSS nfet_03p3 w=0.85u l=0.3u
X24 VSS a_25_21# a_205_70# VSS nfet_03p3 w=0.85u l=0.3u
X25 a_201_111# CLK a_184_21# VDD pfet_03p3 w=1.7u l=0.3u
X26 VSS a_41_111# a_145_21# VSS nfet_03p3 w=0.85u l=0.3u
X27 a_184_21# a_122_16# a_173_111# VDD pfet_03p3 w=1.7u l=0.3u
X28 a_184_21# CLK a_173_21# VSS nfet_03p3 w=0.85u l=0.3u
X29 VDD a_41_111# a_145_111# VDD pfet_03p3 w=1.7u l=0.3u
X30 a_173_111# a_41_111# VDD VDD pfet_03p3 w=1.7u l=0.3u
X31 a_122_16# CLK VSS VSS nfet_03p3 w=0.85u l=0.3u
.ends
