* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffn_1 Q QN D CLK VDD VSS
X0 a_19_16# a_52_83# a_42_111# VDD pfet_03p3 w=1.7u l=0.3u
X1 a_75_111# a_52_16# a_19_16# VDD pfet_03p3 w=1.7u l=0.3u
X2 a_131_21# a_52_16# a_114_21# VSS nfet_03p3 w=0.85u l=0.3u
X3 a_42_111# D VDD VDD pfet_03p3 w=1.7u l=0.3u
X4 VDD a_19_16# a_9_21# VDD pfet_03p3 w=1.7u l=0.3u
X5 VDD a_135_70# QN VDD pfet_03p3 w=1.7u l=0.3u
X6 Q QN VDD VDD pfet_03p3 w=1.7u l=0.3u
X7 a_75_21# a_52_83# a_19_16# VSS nfet_03p3 w=0.85u l=0.3u
X8 VSS a_135_70# a_131_21# VSS nfet_03p3 w=0.85u l=0.3u
X9 Q QN VSS VSS nfet_03p3 w=0.85u l=0.3u
X10 a_19_16# a_52_16# a_42_21# VSS nfet_03p3 w=0.85u l=0.3u
X11 VSS a_19_16# a_9_21# VSS nfet_03p3 w=0.85u l=0.3u
X12 VSS a_135_70# QN VSS nfet_03p3 w=0.85u l=0.3u
X13 a_52_16# a_52_83# VDD VDD pfet_03p3 w=1.7u l=0.3u
X14 VDD a_135_70# a_131_111# VDD pfet_03p3 w=1.7u l=0.3u
X15 VSS CLK a_52_83# VSS nfet_03p3 w=0.85u l=0.3u
X16 a_131_111# a_52_83# a_114_21# VDD pfet_03p3 w=1.7u l=0.3u
X17 a_114_21# a_52_16# a_103_111# VDD pfet_03p3 w=1.7u l=0.3u
X18 a_114_21# a_52_83# a_103_21# VSS nfet_03p3 w=0.85u l=0.3u
X19 a_135_70# a_114_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X20 a_52_16# a_52_83# VSS VSS nfet_03p3 w=0.85u l=0.3u
X21 a_42_21# D VSS VSS nfet_03p3 w=0.85u l=0.3u
X22 VDD a_9_21# a_75_111# VDD pfet_03p3 w=1.7u l=0.3u
X23 a_103_111# a_9_21# VDD VDD pfet_03p3 w=1.7u l=0.3u
X24 a_103_21# a_9_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X25 a_135_70# a_114_21# VSS VSS nfet_03p3 w=0.85u l=0.3u
X26 VSS a_9_21# a_75_21# VSS nfet_03p3 w=0.85u l=0.3u
X27 VDD CLK a_52_83# VDD pfet_03p3 w=1.7u l=0.3u
.ends
