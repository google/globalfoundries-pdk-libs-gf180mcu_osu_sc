# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__tbuf_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__tbuf_1 0 0 ;
  SIZE 5.2 BY 8.3 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 7.6 5.2 8.3 ;
        RECT 3.55 5.55 3.8 8.3 ;
        RECT 1.4 5.55 1.65 8.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 0 5.2 0.7 ;
        RECT 3.55 0 3.8 1.9 ;
        RECT 1.4 0 1.65 1.9 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 4.25 1.55 4.55 ;
      LAYER Metal2 ;
        RECT 1.05 4.25 1.55 4.55 ;
        RECT 1.1 4.2 1.5 4.6 ;
      LAYER Via1 ;
        RECT 1.17 4.27 1.43 4.53 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3 2.35 3.5 2.65 ;
      LAYER Metal2 ;
        RECT 3 2.3 3.5 2.7 ;
      LAYER Via1 ;
        RECT 3.12 2.37 3.38 2.63 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.8 5.55 3.05 7.25 ;
        RECT 1.95 1.65 3.05 1.9 ;
        RECT 2.8 1.05 3.05 1.9 ;
        RECT 2.45 3.6 2.95 3.9 ;
        RECT 1.95 4.35 2.8 4.6 ;
        RECT 2.55 2.85 2.8 4.6 ;
        RECT 1.95 5.55 3.05 5.8 ;
        RECT 1.95 2.85 2.8 3.1 ;
        RECT 1.95 4.35 2.2 5.8 ;
        RECT 1.95 1.65 2.2 3.1 ;
      LAYER Metal2 ;
        RECT 2.45 3.55 2.95 3.95 ;
      LAYER Via1 ;
        RECT 2.57 3.62 2.83 3.88 ;
    END
  END Y
  OBS
    LAYER Metal2 ;
      RECT 4.3 4.85 4.8 5.25 ;
      RECT 2.45 4.85 2.95 5.25 ;
      RECT 2.45 4.9 4.8 5.2 ;
    LAYER Via1 ;
      RECT 4.42 4.92 4.68 5.18 ;
      RECT 2.57 4.92 2.83 5.18 ;
    LAYER Metal1 ;
      RECT 4.4 1.05 4.65 7.25 ;
      RECT 4.3 4.9 4.8 5.2 ;
      RECT 0.55 1.05 0.8 7.25 ;
      RECT 0.55 3.45 2 3.75 ;
      RECT 2.45 4.9 2.95 5.2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__tbuf_1
