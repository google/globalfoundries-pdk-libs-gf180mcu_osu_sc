* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* SKY130 Spice File.
.param sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre = 0.0
.param sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre = 0.0
* statistics {
*   process {
*   }
*   mismatch {
*     vary sky130_fd_pr__pfet_01v8_lvt__toxe_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__vth0_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__voff_slope_spectre dist=gauss std = 1.0
*     vary sky130_fd_pr__pfet_01v8_lvt__nfactor_slope_spectre dist=gauss std = 1.0
*   }
* }
.subckt  sky130_fd_pr__pfet_01v8_lvt d g s b
+ 
.param  l = 1 w = 1 nf = 1.0 ad = 0 as = 0 pd = 0 ps = 0 nrd = 0 nrs = 0 sa = 0 sb = 0 sd = 0 mult = 1

.model sky130_fd_pr__pfet_01v8_lvt.0 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.353895+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.64774
+ k2 = -0.015394
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00239108
+ a0 = 1.75036
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.338792
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.1 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-0.353895+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))}
+ k1 = 0.64774
+ k2 = -0.015394
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.0054e-9
+ ub = 3.0419e-18
+ uc = 4.9353e-11
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 0.00239108
+ a0 = 1.75036
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 0.338792
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 0.0018466
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 0.01363
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.2 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.600368143e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.895115065e-8
+ k1 = 0.64774
+ k2 = -1.748031120e-02 lk2 = 1.662820276e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.063860385e-09 lua = 4.659377462e-16
+ ub = 3.130434233e-18 lub = -7.056306785e-25
+ uc = 3.786240783e-11 luc = 9.158168570e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.311716801e-03 lu0 = 6.325362001e-10
+ a0 = 1.842794901e+00 la0 = -7.367195637e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.220434470e-01 lags = 1.334883956e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 8.564218525e-05 lpdiblc2 = 1.403508912e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.907075439e-03 ldelta = 6.155282858e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112753625e-01 lkt1 = 7.910657830e-8
+ kt2 = -0.055045
+ at = 2.990885676e+05 lat = -1.075058399e-1
+ ute = -3.117702777e-01 lute = 7.098233271e-7
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -1.752002700e-19 lub1 = 2.116892035e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.3 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.180632133e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.176901317e-7
+ k1 = 0.64774
+ k2 = -2.243051758e-02 lk2 = 3.628123989e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.562792134e+05 lvsat = -1.291059924e-1
+ ua = -3.111105615e-09 lua = 6.535081584e-16
+ ub = 3.173159225e-18 lub = -8.752550918e-25
+ uc = 6.007988243e-11 luc = 3.375090010e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.160771715e-03 lu0 = 1.231810082e-9
+ a0 = 2.228193782e+00 la0 = -2.266809005e-6
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.868307461e-01 lags = -1.237265760e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.046519360e-04 lpdiblc2 = 1.316558866e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.970091414e-02 ldelta = 6.789288827e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.767429082e+05 lat = -4.158048318e-1
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.566973875e-19 lub1 = 1.382300769e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.4 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.832630588e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.076301802e-8
+ k1 = 0.64774
+ k2 = 5.917477239e-02 lk2 = -1.244930141e-07 pk2 = 2.524354897e-29
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 90748.0
+ ua = -2.243679162e-09 lua = -1.055447730e-15
+ ub = 1.846518971e-18 lub = 1.738418572e-24
+ uc = 3.314575453e-11 luc = 5.643922743e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.062603080e-03 lu0 = -5.449284742e-10
+ a0 = 1.034947452e+00 la0 = 8.405928658e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.750161028e-01 lags = 2.935789845e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.112108092e-03 lpdiblc2 = 1.989710134e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.706942057e-02 ldelta = 1.197371273e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.051780947e+05 lat = -7.779727233e-2
+ ute = -0.13298
+ ua1 = 7.984120920e-10 lua1 = -2.015893579e-16
+ ub1 = -3.088062225e-19 lub1 = 4.379065378e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.5 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.589178955e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -2.502790205e-8
+ k1 = 0.64774
+ k2 = -4.760978368e-02 lk2 = 3.249576706e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 9.004367473e+04 lvsat = 1.035460274e-3
+ ua = -3.148449927e-09 lua = 2.746964859e-16
+ ub = 3.138238327e-18 lub = -1.605961802e-25
+ uc = 6.942496448e-11 luc = 3.103528315e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.918792644e-03 lu0 = 1.136638720e-9
+ a0 = 9.509980068e-01 la0 = 2.074771433e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.431627920e-03 lags = 5.458330423e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-1.536687805e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -4.150398619e-8
+ nfactor = {2.596284816e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -8.671623232e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 8.369674000e-04 lpdiblc2 = 1.409138775e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.060167601e-02 ldelta = 2.148223505e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.495587000e-01 lkt1 = 8.557522926e-8
+ kt2 = -9.242662714e-02 lkt2 = 5.495641223e-8
+ at = 2.030761951e+05 lat = -7.470717515e-2
+ ute = 5.154157900e-02 lute = -2.712734768e-7
+ ua1 = 6.6129e-10
+ ub1 = -1.051507649e-20 lub1 = -6.246991736e-28
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.6 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.824282744e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -2.219425523e-9
+ k1 = 0.64774
+ k2 = -3.594975770e-03 lk2 = -1.020497876e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 8.270866259e+04 lvsat = 8.151485628e-3
+ ua = -2.793555873e-09 lua = -6.960220609e-17
+ ub = 2.832314703e-18 lub = 1.361940940e-25
+ uc = 7.560659988e-11 luc = -2.893554361e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.080123227e-03 lu0 = 9.979661004e-12
+ a0 = 1.238460259e+00 la0 = -7.140292371e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.025845857e-01 lags = -1.324467039e-7
+ b0 = 2.868730761e-07 lb0 = -2.783084804e-13
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.101312195e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 1.327276669e-8
+ nfactor = {2.478315184e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 2.773141632e-8
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.087771689e-02 lpdiblc2 = 3.515778014e-8
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.192696355e-02 ldelta = 1.049506397e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.949561231e-01 lkt1 = -6.441168771e-8
+ kt2 = -1.675129156e-02 lkt2 = -1.845963620e-8
+ at = 1.888193129e+05 lat = -6.087593212e-2
+ ute = -6.785458400e-02 lute = -1.554418862e-7
+ ua1 = 4.402654326e-10 lua1 = 2.144258789e-16
+ ub1 = 5.417888777e-19 lub1 = -5.364396188e-25 wub1 = -3.214242366e-40 pub1 = -7.663350977e-47
+ uc1 = -2.221711598e-11 luc1 = 1.189020963e-17 puc1 = 1.175494351e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.7 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 7e-06 wmax = 1.0e-4
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.028958654e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 7.403310033e-9
+ k1 = 0.64774
+ k2 = -4.522682480e-02 lk2 = 9.368026901e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.128891965e+05 lvsat = -6.037741502e-3
+ ua = -3.064749110e-09 lua = 5.789793832e-17
+ ub = 3.036628000e-18 lub = 4.013721894e-26
+ uc = 8.292797020e-11 luc = -6.335660010e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.383542224e-03 lu0 = 3.374737368e-10
+ a0 = 1.271386500e+00 la0 = -8.688303098e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.117992250e-01 lags = 4.264579512e-9
+ b0 = -9.562435870e-07 lb0 = 3.061366032e-13
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.845988310e-02 lpdiblc2 = 6.222974768e-08 ppdiblc2 = 5.048709793e-29
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.625998530e-02 ldelta = 8.457915461e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.533030000e-01 lkt1 = 1.003430473e-8
+ kt2 = -0.056015
+ at = 1.321604503e+05 lat = -3.423805119e-2
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.8 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.755847395e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 1.524807771e-7
+ k1 = 0.64774
+ k2 = -1.845732359e-02 wk2 = 2.153543442e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.122852555e-09 wua = 8.257017961e-16
+ ub = 3.233797857e-18 wub = -1.349058823e-24
+ uc = 5.088466180e-11 wuc = -1.076771721e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.427749342e-03 wu0 = -2.577886978e-10
+ a0 = 1.754187897e+00 wa0 = -2.691045254e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.739447700e-01 wags = -2.471270665e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.355393401e-03 wpdiblc2 = -3.576862384e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.393770920e-03 wdelta = 7.196159122e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.9 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.755847395e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 1.524807771e-7
+ k1 = 0.64774
+ k2 = -1.845732359e-02 wk2 = 2.153543442e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.122852555e-09 wua = 8.257017961e-16
+ ub = 3.233797857e-18 wub = -1.349058823e-24
+ uc = 5.088466180e-11 wuc = -1.076771721e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.427749342e-03 wu0 = -2.577886978e-10
+ a0 = 1.754187897e+00 wa0 = -2.691045254e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.739447700e-01 wags = -2.471270665e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.355393401e-03 wpdiblc2 = -3.576862384e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.393770920e-03 wdelta = 7.196159122e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 285600.0
+ ute = -0.22271
+ ua1 = 6.8217e-10
+ ub1 = -1.4864e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.10 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.617339086e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.103931303e-07 wvth0 = 1.193072215e-08 pvth0 = 1.120204318e-12
+ k1 = 0.64774
+ k2 = -8.561527556e-03 lk2 = -7.887092930e-08 wk2 = -6.269983385e-08 pk2 = 6.713673023e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.328343381e-09 lua = 1.637791679e-15 wua = 1.859338734e-15 pua = -8.238236272e-21
+ ub = 3.544999583e-18 lub = -2.480322883e-24 wub = -2.914430892e-24 pub = 1.247624237e-29
+ uc = 1.049472475e-11 luc = 3.219136548e-16 wuc = 1.923972205e-16 puc = -1.619254012e-21
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.177017047e-03 lu0 = 1.998372745e-09 wu0 = 9.469511287e-10 pu0 = -9.601951105e-15
+ a0 = 2.087742736e+00 la0 = -2.658480431e-06 wa0 = -1.722004835e-06 pa0 = 1.351014801e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.127594949e-01 lags = -3.093589859e-07 wags = -6.377417996e-07 pags = 3.113256062e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.137568765e-04 lpdiblc2 = 1.967948574e-08 wpdiblc2 = 1.401792951e-09 ppdiblc2 = -3.968060493e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.199770227e-02 ldelta = 1.226722731e-07 wdelta = 1.258721629e-07 pdelta = -4.296750735e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112753625e-01 lkt1 = 7.910657830e-8
+ kt2 = -0.055045
+ at = 2.990885676e+05 lat = -1.075058399e-1
+ ute = -3.117702777e-01 lute = 7.098233271e-7
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -1.752002700e-19 lub1 = 2.116892035e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.11 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.313755923e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -6.279345480e-07 wvth0 = -6.094216039e-07 pvth0 = 3.587063148e-12
+ k1 = 0.64774
+ k2 = -6.175389152e-02 lk2 = 1.323104685e-07 wk2 = 2.764467792e-07 pk2 = -6.750939279e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 2.380664658e+05 lvsat = -4.538132438e-01 wvsat = -5.749715821e-01 pvsat = 2.282720552e-6
+ ua = -3.641080482e-09 lua = 2.879403318e-15 wua = 3.725769954e-15 pua = -1.564823885e-20
+ ub = 3.989011391e-18 lub = -4.243114140e-24 wub = -5.735512518e-24 pub = 2.367634548e-29
+ uc = 1.067056105e-10 luc = -6.005751222e-17 wuc = -3.277829714e-16 puc = 4.459367757e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.423817442e-03 lu0 = 4.988684391e-09 wu0 = 5.180853390e-09 pu0 = -2.641115700e-14
+ a0 = 3.453231991e+00 la0 = -8.079670772e-06 wa0 = -8.612126414e-06 pa0 = 4.086492975e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 5.535415305e-01 lags = -8.682840807e-07 wags = -1.171991485e-06 pags = 5.234304779e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.424066316e-03 lpdiblc2 = 9.603959680e-09 wpdiblc2 = -1.489966960e-08 ppdiblc2 = 2.503856512e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.341109718e-02 ldelta = -5.760724502e-08 wdelta = -9.638379330e-08 pdelta = 4.527132998e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 5.795015639e+05 lat = -1.220786095e+00 wat = -1.425411192e+00 pat = 5.659089118e-6
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -2.442646491e-19 lub1 = 4.858848026e-25 wub1 = 6.156055547e-25 pub1 = -2.444043315e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.12 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-8.068887603e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 5.059098424e-07 wvth0 = 2.978125961e-06 pvth0 = -3.480925749e-12
+ k1 = 0.64774
+ k2 = 1.799395057e-01 lk2 = -3.438605695e-07 wk2 = -8.489867022e-07 pk2 = 1.542173218e-12
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -3.855277475e+05 lvsat = 7.747577776e-01 wvsat = 3.348260417e+00 pvsat = -5.446615355e-6
+ ua = -5.020595412e-10 lua = -3.304923094e-15 wua = -1.224373920e-14 pua = 1.581400976e-20
+ ub = -7.967233960e-19 lub = 5.185477322e-24 wub = 1.858222645e-23 pub = -2.423312635e-29
+ uc = 7.157120301e-11 luc = 9.162365034e-18 wuc = -2.701342843e-16 puc = 3.323605030e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 6.158272449e-03 lu0 = -4.338878470e-09 wu0 = -2.176282808e-08 pu0 = 2.667180234e-14
+ a0 = -1.079470648e+00 la0 = 8.504106698e-07 wa0 = 1.486454531e-05 pa0 = -5.387517663e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.495020608e-01 lags = -1.057340240e-06 wags = -3.335678040e-06 pags = 9.497081026e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -6.557872667e-03 lpdiblc2 = 2.729968186e-08 wpdiblc2 = 2.422402819e-08 ppdiblc2 = -5.204079247e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.432301148e-03 ldelta = 2.089002699e-08 wdelta = 1.652191718e-07 pdelta = -6.268247391e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.131987617e-01 lkt1 = 4.370742286e-07 wkt1 = 1.559616317e-06 pkt1 = -3.072670289e-12
+ kt2 = -2.056581243e-01 lkt2 = 2.967296938e-07 wkt2 = 1.058823518e-06 pkt2 = -2.086035860e-12
+ at = -8.422733585e+05 lat = 1.580316660e+00 wat = 7.363675892e+00 pat = -1.165668685e-5
+ ute = -0.13298
+ ua1 = 8.444087353e-10 lua1 = -2.922094147e-16 wua1 = -3.233604498e-16 pua1 = 6.370669734e-22
+ ub1 = 4.146282369e-20 lub1 = -7.703974923e-26 wub1 = -2.462422219e-24 pub1 = 3.620117713e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.13 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.998556189e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 5.452660470e-08 wvth0 = 9.908045975e-07 pvth0 = -5.592751832e-13
+ k1 = 0.64774
+ k2 = -1.438858961e-01 lk2 = 1.322097259e-07 wk2 = 6.768295429e-07 pk2 = -7.009979053e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.207959584e+05 lvsat = -4.106549870e-01 wvsat = -2.325217660e+00 pvsat = 2.894220073e-6
+ ua = -3.211673925e-09 lua = 6.786029455e-16 wua = 4.444702731e-16 pua = -2.839497954e-21
+ ub = 3.114441803e-18 lub = -5.645026398e-25 wub = 1.672916572e-25 pub = 2.839497954e-30
+ uc = 1.037031646e-10 luc = -3.807627769e-17 wuc = -2.409787636e-16 puc = 2.894976600e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.778572054e-03 lu0 = 2.099916168e-09 wu0 = 9.857630867e-10 pu0 = -6.771925228e-15
+ a0 = -1.922902058e+00 la0 = 2.090377141e-06 wa0 = 2.020377036e-05 pa0 = -1.323695268e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.518201707e+00 lags = 2.129498616e-06 wags = 1.069721625e-05 pags = -1.113330835e-11
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-8.266602128e-02+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = -1.458883376e-07 wvoff = -4.991556455e-07 pvoff = 7.338311765e-13
+ nfactor = {2.744634224e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -3.048113721e-07 wnfactor = -1.042909390e-06 pnfactor = 1.533228025e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.740781341e-02 lpdiblc2 = -7.933351695e-09 wpdiblc2 = -1.164945057e-07 ppdiblc2 = 1.548358565e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.515940121e-03 ldelta = 3.324379828e-09 wdelta = 3.575317084e-08 pdelta = 1.276513201e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.229065272e-01 lkt1 = 1.573170516e-07 wkt1 = -1.873671200e-07 pkt1 = -5.043513241e-13
+ kt2 = 5.818649717e-02 lkt2 = -9.116015725e-08 wkt2 = -1.058823518e-06 pkt2 = 1.027212342e-12
+ at = 9.264597157e+05 lat = -1.019977426e+00 wat = -5.085449807e+00 pat = 6.645333046e-6
+ ute = 3.339422440e-01 lute = -6.864434024e-07 wute = -1.985301526e-06 pute = 2.918681112e-12
+ ua1 = 5.184758486e-10 lua1 = 1.869591889e-16 wua1 = 1.003996052e-15 pua1 = -1.314339550e-21
+ ub1 = -9.446375166e-21 lub1 = -2.195845082e-27 wub1 = -7.513064355e-27 pub1 = 1.104529400e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.14 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.155743853e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -2.723841269e-08 wvth0 = 2.330200759e-07 pvth0 = 1.758856815e-13
+ k1 = 0.64774
+ k2 = 4.938137267e-03 lk2 = -1.217116602e-08 wk2 = -5.998853557e-08 pk2 = 1.382246942e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.139217128e+04 lvsat = -5.227974994e-02 wvsat = 2.201576898e-01 pvsat = 4.248369040e-7
+ ua = -1.802874549e-09 lua = -6.881367261e-16 wua = -6.964576891e-15 pua = 4.348352106e-21
+ ub = 1.528294728e-18 lub = 9.742900144e-25 wub = 9.167375178e-24 pub = -5.891888073e-30
+ uc = 3.755050077e-11 luc = 2.610139840e-17 wuc = 2.675377257e-16 puc = -2.038370694e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 4.808819158e-03 lu0 = -8.398629091e-10 wu0 = -1.215288452e-08 pu0 = 5.974468054e-15
+ a0 = 9.816365042e-01 la0 = -7.274464232e-07 wa0 = 1.805493600e-06 pa0 = 4.612043533e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.281505911e-01 lags = -4.978883413e-08 wags = -1.797312681e-07 pags = -5.810920983e-13
+ b0 = 4.426471106e-07 lb0 = -4.294318811e-13 wb0 = -1.095105171e-12 pb0 = 1.062410806e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-2.811339787e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))} lvoff = 4.665435892e-08 wvoff = 4.991556455e-07 pvoff = -2.346755310e-13
+ nfactor = {2.329965776e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 9.747714854e-08 wnfactor = 1.042909390e-06 pnfactor = -4.903186352e-13
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -3.920739735e-02 lpdiblc2 = 4.699161195e-08 wpdiblc2 = 1.288592666e-07 ppdiblc2 = -8.319287895e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.195210279e-03 ldelta = 4.605679280e-09 wdelta = 1.246557859e-07 pdelta = 4.140289265e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.147055172e-01 lkt1 = -1.416826174e-07 wkt1 = -1.267177622e-06 pkt1 = 5.432214353e-13
+ kt2 = -1.675129156e-02 lkt2 = -1.845963620e-8
+ at = -2.981473773e+05 lat = 1.680690224e-01 wat = 3.423418685e+00 pat = -1.609503178e-6
+ ute = -3.502552490e-01 lute = -2.267262556e-08 wute = 1.985301526e-06 pute = -9.333795861e-13
+ ua1 = 5.370829407e-10 lua1 = 1.689076116e-16 wua1 = -6.806356019e-16 pua1 = 3.199974250e-22
+ ub1 = 5.407201764e-19 lub1 = -5.359371742e-25 wub1 = 7.513064355e-27 pub1 = -3.532229641e-33
+ uc1 = -2.221711598e-11 luc1 = 1.189020963e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.15 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.0e-06 wmax = 7.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.477187922e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 3.488861952e-08 wvth0 = 1.018117920e-06 pvth0 = -1.932241444e-13
+ k1 = 0.64774
+ k2 = -1.738068242e-02 lk2 = -1.678084532e-09 wk2 = -1.957608314e-07 pk2 = 7.765513543e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -4.267305201e+05 lvsat = 1.725072428e-01 wvsat = 3.793574094e+00 pvsat = -1.255186952e-6
+ ua = -4.083220101e-09 lua = 3.839563338e-16 wua = 7.159940694e-15 pua = -2.292219214e-21
+ ub = 4.536744328e-18 lub = -4.401175230e-25 wub = -1.054594980e-23 pub = 3.376233099e-30
+ uc = 1.569484238e-10 luc = -3.003293813e-17 wuc = -5.203703028e-16 puc = 1.665939506e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.075305232e-03 lu0 = 4.452849958e-10 wu0 = 2.166933178e-09 pu0 = -7.579226378e-16
+ a0 = -3.907199526e+00 la0 = 1.571015392e-06 wa0 = 3.640591548e-05 pa0 = -1.165517181e-11
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.066011333e+00 lags = -2.086323728e-07 wags = -4.599168693e-06 pags = 1.496684310e-12
+ b0 = -1.475490369e-06 lb0 = 4.723708641e-13 wb0 = 3.650350569e-12 pb0 = -1.168641483e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.428236052e-01 lpdiblc2 = 9.570625399e-08 wpdiblc2 = 4.524826305e-07 ppdiblc2 = -2.353427853e-13
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.115481664e-03 ldelta = 5.583453290e-09 wdelta = 1.697379853e-07 pdelta = 2.020772201e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.034830568e-01 lkt1 = -5.915300989e-09 wkt1 = -3.502385850e-07 pkt1 = 1.121271318e-13
+ kt2 = -0.056015
+ at = 1.321604503e+05 lat = -3.423805119e-02 wat = 4.440892099e-16
+ ute = -0.39848
+ ua1 = 8.9635e-10
+ ub1 = -5.9922e-19
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.16 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.462966848e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 5.159284744e-9
+ k1 = 0.64774
+ k2 = -9.199080460e-03 wk2 = -2.503434326e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.110204400e-09 wua = 7.620804644e-16
+ ub = 3.071653080e-18 wub = -5.334563251e-25
+ uc = 3.028167382e-11 wuc = 9.286712539e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.015692271e-03 wu0 = 1.814894626e-9
+ a0 = 1.755663273e+00 wa0 = -3.433172492e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.426940342e-01 wags = -8.993311560e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.302739548e-04 wpdiblc2 = 4.597631442e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.320486445e-02 wdelta = 2.261092738e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899330258e+05 wat = -2.179550128e-2
+ ute = -1.181113622e-01 wute = -5.261403526e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463825844e-19 wub1 = -1.135499892e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.17 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.462966848e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 5.159284744e-9
+ k1 = 0.64774
+ k2 = -9.199080460e-03 wk2 = -2.503434326e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.110204400e-09 wua = 7.620804644e-16
+ ub = 3.071653080e-18 wub = -5.334563251e-25
+ uc = 3.028167382e-11 wuc = 9.286712539e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.015692271e-03 wu0 = 1.814894626e-9
+ a0 = 1.755663273e+00 wa0 = -3.433172492e-8
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.426940342e-01 wags = -8.993311560e-8
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 7.302739548e-04 wpdiblc2 = 4.597631442e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.320486445e-02 wdelta = 2.261092738e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.60135
+ kt2 = -0.055045
+ at = 2.899330258e+05 wat = -2.179550128e-2
+ ute = -1.181113622e-01 wute = -5.261403526e-7
+ ua1 = 6.8217e-10
+ ub1 = -1.463825844e-19 wub1 = -1.135499892e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.18 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.468345485e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 4.286852149e-09 wvth0 = -6.301437005e-08 pvth0 = 5.433539139e-13
+ k1 = 0.64774
+ k2 = -1.456387440e-02 lk2 = 4.275818560e-08 wk2 = -3.250750102e-08 pk2 = 5.956215099e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.155316483e-09 lua = 3.595498405e-16 wua = 9.889982103e-16 pua = -1.808567338e-21
+ ub = 3.071653080e-18 wub = -5.334563251e-25
+ uc = 3.028167382e-11 wuc = 9.286712539e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.813807988e-03 lu0 = 1.609047016e-09 wu0 = 2.773924659e-09 pu0 = -7.643608426e-15
+ a0 = 1.828132703e+00 la0 = -5.775918641e-07 wa0 = -4.161435242e-07 pa0 = 3.043095403e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.845346156e-01 lags = 4.635389995e-07 wags = 7.240627115e-09 pags = -7.744888197e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.508788799e-03 lpdiblc2 = 1.784565481e-08 wpdiblc2 = 8.418926283e-09 ppdiblc2 = -3.045627397e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.180915593e-02 ldelta = 1.112399932e-08 wdelta = 6.121571177e-09 pdelta = 1.314225599e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.112753625e-01 lkt1 = 7.910657830e-8
+ kt2 = -0.055045
+ at = 3.077222787e+05 lat = -1.417829247e-01 wat = -4.342832639e-02 pat = 1.724167529e-7
+ ute = -1.033537003e-01 lute = -1.176207057e-07 wute = -1.048353725e-06 pute = 4.162116300e-12
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -1.707022877e-19 lub1 = 1.938315615e-25 wub1 = -2.262524697e-26 pub1 = 8.982551111e-32
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.19 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.889279480e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 1.714037516e-07 wvth0 = 1.830806100e-07 pvth0 = -4.336788407e-13
+ k1 = 0.64774
+ k2 = -6.882102049e-03 lk2 = 1.226043551e-08 wk2 = 4.368494803e-10 pk2 = -7.123169742e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.918085040e-09 lua = -5.822933868e-16 wua = 8.903925618e-17 pua = 1.764400204e-21
+ ub = 2.777821499e-18 lub = 1.166553981e-24 wub = 3.568792217e-25 pub = -3.534761219e-30
+ uc = -2.383493495e-12 luc = 1.296854507e-16 wuc = 2.209448215e-16 puc = -5.084870250e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.361054375e-03 lu0 = -5.636004928e-10 wu0 = 4.664691400e-10 pu0 = 1.517324567e-15
+ a0 = 1.336338188e+00 la0 = 1.374903671e-06 wa0 = 2.036035704e-06 pa0 = -6.692411699e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.047720002e-01 lags = 3.831936483e-07 wags = 7.934114444e-08 pags = -1.060738328e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.426316039e-03 lpdiblc2 = 1.751822599e-08 wpdiblc2 = 4.468092478e-09 ppdiblc2 = -1.477089090e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.266170667e-02 ldelta = 7.739249232e-09 wdelta = 7.987466914e-09 pdelta = 1.240146833e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 2.850358334e+05 lat = -5.171444741e-02 wat = 5.577734496e-02 pat = -2.214441472e-7
+ ute = -0.13298
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.20 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.525445780e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -2.943057630e-07 wvth0 = -3.132828588e-07 pvth0 = 5.442291656e-13
+ k1 = 0.64774
+ k2 = 1.372843900e-02 lk2 = -2.834531888e-08 wk2 = -1.293041029e-08 pk2 = -4.489625742e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 5.170091150e+05 lvsat = -7.747577776e-01 wvsat = -1.191579424e+00 pvsat = 2.347584245e-6
+ ua = -3.008063832e-09 lua = -4.050221185e-16 wua = 3.616829159e-16 pua = 1.227252661e-21
+ ub = 2.900357420e-18 lub = 9.251404505e-25 wub = -1.441539975e-26 pub = -2.803256977e-30
+ uc = -3.260388439e-11 luc = 1.892240027e-16 wuc = 2.538755728e-16 puc = -5.733653799e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.084834834e-03 lu0 = 1.950737055e-09 wu0 = 3.757009587e-09 pu0 = -4.965517241e-15
+ a0 = 1.931906820e+00 la0 = 2.015471091e-07 wa0 = -2.829483537e-07 pa0 = -2.123676853e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -3.263049289e-01 lags = 1.626506705e-06 wags = 1.572716990e-06 pags = -4.002905283e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.264540780e-03 lpdiblc2 = 2.902037528e-08 wpdiblc2 = 2.777863099e-08 ppdiblc2 = -6.069603178e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.450525721e-02 ldelta = 6.126210730e-08 wdelta = 2.058268513e-07 pdelta = -2.657575906e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -3.695012383e-01 lkt1 = -4.370742286e-07 wkt1 = -6.722212706e-07 pkt1 = 1.324373375e-12
+ kt2 = 9.556812431e-02 lkt2 = -2.967296938e-07 wkt2 = -4.563710206e-07 pkt2 = 8.991170844e-13
+ at = 1.103455934e+06 lat = -1.664120716e+00 wat = -2.423513672e+00 pat = 4.663118654e-6
+ ute = -0.13298
+ ua1 = 9.074379203e-10 lua1 = -4.163860484e-16 wua1 = -6.404027971e-16 pua1 = 1.261686369e-21
+ ub1 = -9.422767207e-19 lub1 = 1.616300497e-24 wub1 = 2.485874259e-24 pub1 = -4.897532741e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.21 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.213155640e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -4.618794177e-08 wvth0 = 9.273240991e-08 pvth0 = -5.267215164e-14
+ k1 = 0.64774
+ k2 = 6.599456522e-02 lk2 = -1.051841030e-07 wk2 = -3.788876472e-07 pk2 = 4.931139447e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -2.917903252e+05 lvsat = 4.142946754e-01 wvsat = 1.259154054e+00 pvsat = -1.255349324e-6
+ ua = -3.165100539e-09 lua = -1.741553893e-16 wua = 2.102020406e-16 pua = 1.449951512e-21
+ ub = 3.635763045e-18 lub = -1.560124526e-25 wub = -2.455000065e-24 pub = 7.847563658e-31
+ uc = 1.588276526e-10 luc = -9.220811420e-17 wuc = -5.182597888e-16 puc = 5.617855613e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.265889856e-03 lu0 = -1.255730081e-09 wu0 = -6.495576343e-09 pu0 = 1.010727070e-14
+ a0 = 2.527787657e+00 la0 = -6.744841242e-07 wa0 = -2.183590567e-06 pa0 = 6.705427939e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.087696345e+00 lags = -4.522801982e-07 wags = -2.410680273e-06 pags = 1.853266286e-12
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {6.732732404e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = -6.167893972e-06 wnfactor = -2.110339419e-05 pnfactor = 3.102504945e-11
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.429758913e-02 lpdiblc2 = 3.935997614e-08 wpdiblc2 = 4.298645917e-08 ppdiblc2 = -8.305374436e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.786461912e-02 ldelta = -1.572920455e-08 wdelta = -1.269635312e-07 pdelta = 2.234925262e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.525883561e-01 lkt1 = 2.731338822e-07 wkt1 = 9.679526914e-07 pkt1 = -1.086920174e-12
+ kt2 = -2.430397514e-01 lkt2 = 2.010729817e-07 wkt2 = 4.563710206e-07 pkt2 = -4.427460638e-13
+ at = -6.389331553e+05 lat = 8.974438914e-01 wat = 2.788614088e+00 pat = -2.999464913e-6
+ ute = -6.651004501e-01 lute = 7.822942190e-07 wute = 3.039971141e-06 pute = -4.469198373e-12
+ ua1 = 5.907595253e-10 lua1 = 4.917711057e-17 wua1 = 6.404027971e-16 pua1 = -6.212835716e-22
+ ub1 = 4.832609481e-19 lub1 = -4.794465788e-25 wub1 = -2.485874259e-24 pub1 = 2.411658483e-30
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.22 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.628617479e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -5.882119210e-09 wvth0 = -3.212912887e-08 pvth0 = 6.846164590e-14
+ k1 = 0.64774
+ k2 = -5.498372186e-02 lk2 = 1.218237730e-08 wk2 = 2.414236890e-07 pk2 = -1.086779966e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.235512840e+04 lvsat = 9.982658430e-02 wvsat = 3.159156907e-01 pvsat = -3.402713426e-7
+ ua = -3.844482275e-09 lua = 4.849434051e-16 wua = 3.304889636e-15 pua = -1.552344184e-21
+ ub = 3.985761580e-18 lub = -4.955617816e-25 wub = -3.193899345e-24 pub = 1.501595808e-30
+ uc = 7.397815817e-11 luc = -9.891801462e-18 wuc = 8.430340331e-17 puc = -2.278810675e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 7.499305010e-04 lu0 = 1.185115308e-09 wu0 = 8.263682609e-09 pu0 = -4.211350575e-15
+ a0 = 1.685797894e+00 la0 = 1.423680343e-07 wa0 = -1.736500157e-06 pa0 = 2.368002685e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 8.357172459e-01 lags = -2.078239349e-07 wags = -7.208010073e-07 pags = 2.138383659e-13
+ b0 = -2.583528364e-07 lb0 = 2.506397125e-13 wb0 = 2.430986251e-12 pb0 = -2.358409156e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {3.750292032e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 1.087641239e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -7.956673939e-03 lpdiblc2 = 3.320836898e-08 wpdiblc2 = -2.833462217e-08 ppdiblc2 = -1.386195389e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.507652752e-03 ldelta = 1.760203459e-08 wdelta = 1.281142608e-07 pdelta = -2.396991826e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.363242103e-01 lkt1 = -3.368819752e-08 wkt1 = -1.524160929e-07 pkt1 = -8.077935669e-28
+ kt2 = -9.569980137e-03 lkt2 = -2.542654958e-08 wkt2 = -3.612262842e-08 pkt2 = 3.504418734e-14
+ at = 5.044506308e+05 lat = -2.118041718e-01 wat = -6.137199244e-01 pat = 3.012924181e-7
+ ute = 5.977019803e-01 lute = -4.428072448e-07 wute = -2.783006758e-06 pute = 1.179934521e-12
+ ua1 = 4.017700790e-10 lua1 = 2.325242770e-16
+ ub1 = 4.910001242e-19 lub1 = -4.869547018e-25 wub1 = 2.576093020e-25 pub1 = -2.499183763e-31
+ uc1 = -2.221711598e-11 luc1 = 1.189020963e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.23 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 3.0e-06 wmax = 5.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.641879554e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -5.227310937e-08 wvth0 = -4.080671400e-07 pvth0 = 2.452070221e-13
+ k1 = 0.64774
+ k2 = -1.982450596e-02 lk2 = -4.347552259e-09 wk2 = -1.834681839e-07 pk2 = 9.108279301e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 6.571067022e+05 lvsat = -1.938972444e-01 wvsat = -1.658222511e+00 pvsat = 5.878598624e-7
+ ua = -2.881902319e-09 lua = 3.239125145e-17 wua = 1.117206531e-15 pua = -5.238159114e-22
+ ub = 2.744771912e-18 lub = 8.788330586e-26 wub = -1.532170852e-24 pub = 7.203424651e-31
+ uc = -9.645009569e-12 luc = 2.942321273e-17 wuc = 3.176093274e-16 puc = -1.324757204e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.573962792e-03 lu0 = 7.977006465e-10 wu0 = 4.688729771e-09 pu0 = -2.530604373e-15
+ a0 = 5.695994422e+00 la0 = -1.743005812e-06 wa0 = -1.189899516e-05 pa0 = 5.014646483e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -8.197089804e-02 lags = 2.236225575e-07 wags = 1.175282954e-06 pags = -6.775960279e-13
+ b0 = 8.611761213e-07 lb0 = -2.757012294e-13 wb0 = -8.103287502e-12 pb0 = 2.594226977e-18
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {3.750292032e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = 1.087641239e-5
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -2.396427630e-02 lpdiblc2 = 4.073426319e-08 wpdiblc2 = -1.453902536e-07 ppdiblc2 = 4.117116594e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.829745305e-02 ldelta = -8.157116069e-09 wdelta = -1.128622748e-07 pdelta = 8.932399506e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.751464801e-01 lkt1 = 3.157839851e-08 wkt1 = 1.023474064e-08 pkt1 = -7.646947612e-14
+ kt2 = -7.995270474e-02 lkt2 = 7.663536486e-09 wkt2 = 1.204087614e-07 pkt2 = -3.854826291e-14
+ at = 1.152554257e+05 lat = -2.882599209e-02 wat = 8.503376126e-02 pat = -2.722313350e-8
+ ute = -2.281951176e-01 lute = -5.451585367e-08 wute = -8.565479435e-07 pute = 2.742195414e-13
+ ua1 = 8.9635e-10
+ ub1 = -4.285077434e-19 lub1 = -5.465267539e-26 wub1 = -8.586976734e-25 pub1 = 2.749077667e-31
+ uc1 = 3.0734e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.24 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.576745725e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 3.963528567e-8
+ k1 = 0.64774
+ k2 = -2.442027453e-02 wk2 = 2.108721424e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844484786e-09 wua = -4.307335057e-17
+ ub = 2.872732046e-18 wub = 6.929191179e-26
+ uc = 5.904699914e-11 wuc = 5.705658322e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.625531850e-03 wu0 = -3.297296199e-11
+ a0 = 1.865421390e+00 wa0 = -3.669084761e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.939442028e-01 wags = -2.452256364e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.688168638e-03 wpdiblc2 = -1.334961742e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.466374144e-02 wdelta = -1.211047828e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.910491200e-01 wkt1 = -3.121257288e-8
+ kt2 = -0.055045
+ at = 2.871075731e+05 wat = -1.323413090e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.25 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.576745725e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 3.963528567e-8
+ k1 = 0.64774
+ k2 = -2.442027453e-02 wk2 = 2.108721424e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.844484786e-09 wua = -4.307335057e-17
+ ub = 2.872732046e-18 wub = 6.929191179e-26
+ uc = 5.904699914e-11 wuc = 5.705658322e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.625531850e-03 wu0 = -3.297296199e-11
+ a0 = 1.865421390e+00 wa0 = -3.669084761e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.939442028e-01 wags = -2.452256364e-7
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.688168638e-03 wpdiblc2 = -1.334961742e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.466374144e-02 wdelta = -1.211047828e-8
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.910491200e-01 wkt1 = -3.121257288e-8
+ kt2 = -0.055045
+ at = 2.871075731e+05 wat = -1.323413090e-2
+ ute = -0.29175
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.26 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.884345460e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 2.451614494e-07 wvth0 = 6.303728309e-08 pvth0 = -1.865173127e-13
+ k1 = 0.64774
+ k2 = -3.812456051e-02 lk2 = 1.092251464e-07 wk2 = 3.888345122e-08 pk2 = -1.418385892e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.824932695e-09 lua = -1.558329979e-16 wua = -1.209374053e-17 pua = -2.469119840e-22
+ ub = 2.915161633e-18 lub = -3.381699587e-25 wub = -5.927346986e-26 pub = 1.024684734e-30
+ uc = 5.904699914e-11 wuc = 5.705658322e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.807751003e-03 lu0 = -1.452313071e-09 wu0 = -2.378101435e-10 pu0 = 1.632582038e-15
+ a0 = 1.828620667e+00 la0 = 2.933070948e-07 wa0 = -4.176220977e-07 pa0 = 4.041949179e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.843327173e-01 lags = 7.660493305e-08 wags = -2.951564033e-07 pags = 3.979554520e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.835833599e-03 lpdiblc2 = -1.176911153e-09 wpdiblc2 = -4.745661909e-09 ppdiblc2 = 2.718377488e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.928614596e-02 ldelta = 4.286021574e-08 wdelta = -1.653436659e-08 pdelta = 3.525903132e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.907504857e-01 lkt1 = -2.380158728e-09 wkt1 = -6.219218291e-08 pkt1 = 2.469119840e-13
+ kt2 = -0.055045
+ at = 3.020924617e+05 lat = -1.194317350e-01 wat = -2.636948556e-02 pat = 1.046906812e-7
+ ute = -4.493349804e-01 lute = 1.255975144e-06 pute = -4.038967835e-28
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -1.526239818e-19 lub1 = 1.987739690e-26 wub1 = -7.740410466e-26 pub1 = 6.169219377e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.27 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.408083627e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 5.607859587e-08 wvth0 = 3.727403201e-08 pvth0 = -8.423347030e-14
+ k1 = 0.64774
+ k2 = -8.354699488e-03 lk2 = -8.965518503e-09 wk2 = 4.898949310e-09 pk2 = -6.915188888e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.838816122e-09 lua = -1.007137809e-16 wua = -1.511525414e-16 pua = 3.051716191e-22
+ ub = 2.799288376e-18 lub = 1.218636749e-25 wub = 2.918326970e-25 pub = -3.692576591e-31
+ uc = 7.359668147e-11 luc = -5.776434857e-17 wuc = -9.281794854e-18 puc = 5.950236229e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.518422352e-03 lu0 = -3.036363740e-10 wu0 = -1.036967774e-11 pu0 = 7.296104103e-16
+ a0 = 2.161710405e+00 la0 = -1.029107465e-06 wa0 = -4.649147478e-07 pa0 = 5.919535964e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.395141476e-01 lags = -1.424733464e-07 wags = -3.289394195e-07 pags = 5.320789247e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.790679280e-05 lpdiblc2 = 9.931263967e-09 wpdiblc2 = 3.136844652e-11 ppdiblc2 = 8.218271702e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.222232687e-02 ldelta = 7.090460177e-08 wdelta = 9.318826383e-09 pdelta = -6.738189349e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.034436635e+05 lat = -1.247962019e-1
+ ute = -1.437765289e-01 lute = 4.286378517e-08 wute = 3.271443262e-08 pute = -1.298810411e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.729703344e-19 lub1 = 1.006553670e-25 wub1 = 1.548082093e-25 pub1 = -3.049946195e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.28 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.241417248e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.737715976e-07 wvth0 = -9.633720354e-08 pvth0 = 1.790000374e-13
+ k1 = 0.64774
+ k2 = 2.028634749e-02 lk2 = -6.539253401e-08 wk2 = -3.280145013e-08 pk2 = 6.736006457e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.889936106e-09 wua = 3.745508745e-18
+ ub = 2.861143556e-18 wub = 1.044060563e-25
+ uc = 4.427683518e-11 wuc = 2.092022697e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.124375099e-03 lu0 = 4.726938507e-10 wu0 = 6.071111034e-10 pu0 = -4.869162633e-16
+ a0 = 2.023333902e+00 la0 = -7.564856880e-07 wa0 = -5.599804577e-07 pa0 = 7.792468294e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.323032930e-01 lags = 4.627765828e-07 wags = 1.830937199e-07 pags = -4.767006046e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.833968416e-03 lpdiblc2 = 1.361912955e-08 wpdiblc2 = 1.132351883e-08 ppdiblc2 = -1.402890192e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 6.854742426e-02 ldelta = -4.006400721e-08 wdelta = -4.583008223e-08 pdelta = 4.126945306e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -0.59135
+ kt2 = -0.055045
+ at = 3.363653911e+05 lat = -1.896567789e-01 wat = -9.916182419e-02 pat = 1.953631721e-7
+ ute = -1.220198637e-01 wute = -3.321017754e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.29 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-2.322042681e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = -1.619184898e-07 wvth0 = -1.772826585e-07 pvth0 = 2.980015933e-13
+ k1 = 0.64774
+ k2 = -6.225593716e-02 lk2 = 5.595659306e-08 wk2 = 9.722661018e-09 pk2 = 4.843455185e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.203594064e-09 lua = 4.611226785e-16 wua = 3.268408073e-16 pua = -4.749969377e-22
+ ub = 2.755023104e-18 lub = 1.560124526e-25 wub = 2.137194609e-25 pub = -1.607065553e-31
+ uc = -5.176364414e-11 luc = 1.411934305e-16 wuc = 1.198503722e-16 puc = -1.454416584e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.569897409e-04 lu0 = 3.218021098e-09 wu0 = 2.621655789e-09 pu0 = -3.448589060e-15
+ a0 = 1.940412040e+00 la0 = -6.345785269e-07 wa0 = -4.037907575e-07 pa0 = 5.496253225e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.877485659e-01 lags = 2.342494920e-07 wags = 1.323189332e-08 pags = -2.269790896e-13
+ b0 = 0.0
+ b1 = 2.1073e-24
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {-1.658132404e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} lnfactor = 6.167893972e-06 wnfactor = 4.321664575e-06 pnfactor = -6.353473566e-12
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 3.718040469e-03 lpdiblc2 = 5.456871448e-09 wpdiblc2 = -1.160248389e-08 ppdiblc2 = 1.967564635e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 4.180797482e-03 ldelta = 5.456426730e-08 wdelta = -2.489858747e-08 pdelta = 1.049712070e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.290640143e-01 lkt1 = -9.156943040e-08 wkt1 = -1.235453438e-08 pkt1 = 1.816295694e-14
+ kt2 = -9.242662714e-02 lkt2 = 5.495641223e-8
+ at = 2.269934913e+05 lat = -2.886422726e-02 wat = 1.647801477e-01 pat = -1.926697982e-7
+ ute = 5.871928651e-01 lute = -1.042645547e-06 wute = -7.545878062e-07 pute = 1.060529714e-12
+ ua1 = 8.021074456e-10 lua1 = -1.558610176e-16
+ ub1 = -3.371357726e-19 lub1 = 3.164571978e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.30 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-4.024858381e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 3.279323940e-09 wvth0 = 8.793535152e-08 pvth0 = 4.070166694e-14
+ k1 = 0.64774
+ k2 = 2.987184033e-02 lk2 = -3.342070963e-08 wk2 = -1.569613177e-08 pk2 = 2.950336991e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.311964600e+05 lvsat = -7.214444471e-03 wvsat = 1.641775796e-02 pvsat = -1.592760580e-8
+ ua = -2.704915118e-09 lua = -2.266820703e-17 wua = -1.480991325e-16 pua = -1.423632982e-23
+ ub = 2.954579903e-18 lub = -3.758657786e-26 wub = -6.932811837e-26 pub = 1.138906385e-31
+ uc = 1.172139814e-10 luc = -2.273936810e-17 wuc = -4.670494594e-17 puc = 1.614115075e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.822208051e-03 lu0 = -2.407576196e-10 wu0 = -1.045588728e-09 pu0 = 1.091698716e-16
+ a0 = 8.055535892e-01 la0 = 4.663987244e-07 wa0 = 9.307175478e-07 pa0 = -7.450412373e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.154787499e-01 lags = -1.807108074e-07 wags = -3.564677837e-07 pags = 1.316832035e-13
+ b0 = 9.038980076e-07 lb0 = -8.769121326e-13 wb0 = -1.090736085e-12 pb0 = 1.058172159e-18
+ b1 = 1.599951261e-07 lb1 = -1.552184716e-13 wb1 = -4.847993116e-13 pb1 = 4.703256281e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {4.699570797e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -2.227329201e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.998401769e-02 lpdiblc2 = 2.845130466e-08 wpdiblc2 = 8.109287808e-09 ppdiblc2 = 5.523695969e-16
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 5.259014897e-02 ldelta = 7.600177004e-09 wdelta = -2.061002205e-08 pdelta = 6.336590401e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.810165615e-01 lkt1 = -4.116792651e-08 wkt1 = -1.699433577e-08 pkt1 = 2.266423707e-14
+ kt2 = -2.149129345e-02 lkt2 = -1.386114707e-8
+ at = 3.225041544e+05 lat = -1.215234196e-01 wat = -6.240608968e-02 pat = 2.773379412e-8
+ ute = -4.407998051e-01 lute = -4.534359814e-08 wute = 3.637450404e-07 pute = -2.441530563e-14
+ ua1 = 4.017700790e-10 lua1 = 2.325242770e-16
+ ub1 = 5.760172267e-19 lub1 = -5.694336187e-25 wub1 = -9.183549616e-41 pub1 = -5.473822126e-48
+ uc1 = -2.221711598e-11 luc1 = 1.189020963e-17
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.31 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 1e-06 wmax = 3.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.139074115e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} lvth0 = 5.566361955e-08 wvth0 = 3.486047872e-07 pvth0 = -8.185076490e-14
+ k1 = 0.64774
+ k2 = -1.035080946e-01 lk2 = 2.928719988e-08 wk2 = 7.010045382e-08 pk2 = -1.083346582e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.049218478e+05 lvsat = 5.138433080e-03 wvsat = 1.494618978e-02 pvsat = -1.523575537e-8
+ ua = -2.344402630e-09 lua = -1.921613508e-16 wua = -5.114648255e-16 pua = 1.565982339e-22
+ ub = 2.070038343e-18 lub = 3.782762137e-25 wub = 5.123312397e-25 pub = -1.595736004e-31
+ uc = 1.149190090e-10 luc = -2.166039830e-17 wuc = -5.983061062e-17 puc = 2.231211637e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.690227517e-03 lu0 = -1.787076316e-10 wu0 = -1.723738578e-09 pu0 = 4.279986331e-16
+ a0 = 2.081342933e+00 la0 = -1.334072566e-07 wa0 = -9.462830616e-07 pa0 = 1.374212142e-13
+ keta = -1.175005990e-02 lketa = -3.901921878e-10 wketa = -2.514791535e-09 pketa = 1.182316666e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.311062534e-01 wags = -7.637716583e-8
+ b0 = -3.019344434e-06 lb0 = 9.675806852e-13 wb0 = 3.655031266e-12 pb0 = -1.173026632e-18
+ b1 = -3.086506533e-07 lb1 = 6.511299834e-14 wb1 = 9.352386406e-13 pb1 = -1.972981149e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {4.699570797e+00+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))} wnfactor = -2.227329201e-6
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -8.768161324e-02 lpdiblc2 = 6.027899072e-08 wpdiblc2 = 4.767888446e-08 ppdiblc2 = -1.805107842e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -1.082909500e-02 ldelta = 3.741641746e-08 wdelta = 9.659724891e-08 pdelta = -4.876782200e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.772329190e-01 lkt1 = 4.067712875e-09 wkt1 = 1.655683413e-08 pkt1 = 6.890322292e-15
+ kt2 = -7.244964729e-02 lkt2 = 1.009666820e-08 wkt2 = 9.767383703e-08 pkt2 = -4.592086611e-14
+ at = 1.450285966e+05 lat = -3.808417342e-02 wat = -5.181566450e-03 pat = 8.299706397e-10
+ ute = -6.288086517e-01 lute = 4.304782103e-08 wute = 3.573463186e-07 pute = -2.140697858e-14
+ ua1 = 7.059804287e-10 lua1 = 8.950130210e-17 wua1 = 5.768365536e-16 pua1 = -2.711968215e-22
+ ub1 = -3.087450634e-19 lub1 = -1.534670518e-25 wub1 = -1.221589133e-24 pub1 = 5.743240229e-31
+ uc1 = 3.267269148e-11 luc1 = -1.391595889e-17 wuc1 = -8.968845793e-17 puc1 = 4.216658005e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.32 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.410637394e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope/sqrt(1))} wvth0 = 2.252466589e-8
+ k1 = 0.64774
+ k2 = -5.865868569e-03 wk2 = 1.974543310e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.700285115e-09 wua = -1.916117012e-16
+ ub = 2.763395431e-18 wub = 1.819182472e-25
+ uc = 7.041395077e-11 wuc = -6.003302156e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.109242146e-03 wu0 = -5.312371342e-10
+ a0 = 1.232502242e+00 wa0 = 2.850539425e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.572105307e-02 wags = 1.443774914e-7
+ b0 = -7.512139600e-08 wb0 = 7.738164856e-14
+ b1 = -2.786098210e-07 wb1 = 2.869926333e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.628792926e-03 wpdiblc2 = -1.273799534e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.204718068e-02 wdelta = 8.856895683e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.527707076e-01 wkt1 = -7.064270620e-8
+ kt2 = -0.055045
+ at = 2.640117787e+05 wat = 1.055656982e-2
+ ute = -2.992653623e-01 wute = 7.741484532e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.33 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.410637394e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} wvth0 = 2.252466589e-8
+ k1 = 0.64774
+ k2 = -5.865868569e-03 wk2 = 1.974543310e-9
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.700285115e-09 wua = -1.916117012e-16
+ ub = 2.763395431e-18 wub = 1.819182472e-25
+ uc = 7.041395077e-11 wuc = -6.003302156e-18
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.109242146e-03 wu0 = -5.312371342e-10
+ a0 = 1.232502242e+00 wa0 = 2.850539425e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.572105307e-02 wags = 1.443774914e-7
+ b0 = -7.512139600e-08 wb0 = 7.738164856e-14
+ b1 = -2.786098210e-07 wb1 = 2.869926333e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.628792926e-03 wpdiblc2 = -1.273799534e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.204718068e-02 wdelta = 8.856895683e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.527707076e-01 wkt1 = -7.064270620e-8
+ kt2 = -0.055045
+ at = 2.640117787e+05 wat = 1.055656982e-2
+ ute = -2.992653623e-01 wute = 7.741484532e-9
+ ua1 = 6.8217e-10
+ ub1 = -1.5013e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.34 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.221060390e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -1.510956209e-07 wvth0 = -5.286915996e-09 pvth0 = 2.216623403e-13
+ k1 = 0.64774
+ k2 = 1.846939561e-02 lk2 = -1.939555842e-07 wk2 = -1.941330385e-08 pk2 = 1.704642431e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.638247511e-09 lua = -4.944486993e-16 wua = -2.043959086e-16 pua = 1.018919866e-22
+ ub = 2.614226952e-18 lub = 1.188894411e-24 wub = 2.507157343e-25 pub = -5.483259484e-31
+ uc = 6.349717358e-11 luc = 5.512771719e-17 wuc = 1.121587033e-18 puc = -5.678639994e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.978028765e-03 lu0 = 1.045789678e-09 wu0 = -4.132112229e-10 pu0 = -9.406836270e-16
+ a0 = 9.914238689e-01 la0 = 1.921429592e-06 wa0 = 4.447642776e-07 pa0 = -1.272914529e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -1.510923007e-01 lags = 1.329526617e-06 wags = 2.563784826e-07 pags = -8.926641397e-13
+ b0 = -2.356543279e-08 lb0 = -4.109085024e-13 wb0 = 2.427446953e-14 pb0 = 4.232719174e-19
+ b1 = -3.018064859e-07 lb1 = 1.848807830e-13 wb1 = 3.108872394e-13 pb1 = -1.904434759e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = -1.229392630e-03 lpdiblc2 = 3.075029832e-08 wpdiblc2 = -5.581211529e-10 ppdiblc2 = -5.704060469e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -4.362737452e-03 ldelta = 1.307894269e-07 wdelta = 7.826064424e-09 pdelta = -5.531579395e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.825723843e-01 lkt1 = 2.375236850e-07 wkt1 = -7.061634701e-08 pkt1 = -2.100865703e-16
+ kt2 = -0.055045
+ at = 2.525547307e+05 lat = 9.131433359e-02 wat = 2.465873673e-02 pat = -1.123963151e-7
+ ute = -4.166700854e-01 lute = 9.357326667e-07 wute = -3.364771637e-08 pute = 3.298779326e-13
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -2.917032256e-19 lub1 = 1.128359136e-24 wub1 = 6.585975539e-26 pub1 = -5.249118001e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.35 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.322076224e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -1.109908703e-07 wvth0 = 2.841451263e-08 pvth0 = 8.786278192e-14
+ k1 = 0.64774
+ k2 = -2.598164182e-02 lk2 = -1.747852015e-08 wk2 = 2.305625108e-08 pk2 = 1.853951956e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.888233357e-09 lua = 4.980313584e-16 wua = -1.002484403e-16 pua = -3.115885641e-22
+ ub = 3.075504777e-18 lub = -6.424454416e-25 wub = 7.305496539e-27 pub = 4.180479901e-31
+ uc = 7.738274128e-11 wuc = -1.318176963e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.053280854e-03 lu0 = 7.470279706e-10 wu0 = -5.613210032e-10 pu0 = -3.526663231e-16
+ a0 = 1.737414518e+00 la0 = -1.040261453e-06 wa0 = -2.785264568e-08 pa0 = 6.034431857e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.093212751e-02 lags = 4.480574438e-07 wags = 5.073249643e-08 pags = -7.621975591e-14
+ b0 = -1.810815772e-07 lb0 = 2.144534308e-13 wb0 = 1.865299597e-13 pb0 = -2.209059056e-19
+ b1 = -2.578038001e-07 lb1 = 1.018373996e-14 wb1 = 2.655606008e-13 pb1 = -1.049014832e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.376759897e-03 lpdiblc2 = 2.040349489e-08 wpdiblc2 = -1.347768070e-09 ppdiblc2 = -2.569047711e-15
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.366730071e-02 ldelta = -2.019533894e-08 wdelta = -1.277138383e-08 pdelta = 2.645906223e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.227449259e-01 wkt1 = -7.066926360e-8
+ kt2 = -0.055045
+ at = 3.003473739e+05 lat = -9.842939001e-02 wat = 3.189450696e-03 pat = -2.716013650e-8
+ ute = -1.329931974e-01 lute = -1.905057119e-07 wute = 2.160665223e-08 pute = 1.105100774e-13
+ ua1 = 6.9609e-10
+ ub1 = 1.051881531e-19 lub1 = -4.473571865e-25 wub1 = -1.317195108e-25 pub1 = 2.595065356e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.36 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.885440191e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} wvth0 = 7.301162702e-8
+ k1 = 0.64774
+ k2 = -3.485333408e-02 wk2 = 2.399727418e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -2.635444167e-09 wua = -2.584035832e-16
+ ub = 2.749414341e-18 wub = 2.194969800e-25
+ uc = 7.738274128e-11 wuc = -1.318176963e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 3.432454961e-03 wu0 = -7.403262658e-10
+ a0 = 1.209401883e+00 wa0 = 2.784411478e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.983557150e-01 wags = 1.204511255e-8
+ b0 = -7.222997959e-08 wb0 = 7.440323522e-14
+ b1 = -2.526347694e-07 wb1 = 2.602360444e-13
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.173310164e-02 wpdiblc2 = -2.651757223e-9
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.341661412e-02 wdelta = 6.586237269e-10
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -5.227449259e-01 wkt1 = -7.066926360e-8
+ kt2 = -0.055045
+ at = 2.503868939e+05 wat = -1.059640593e-2
+ ute = -2.296894872e-01 wute = 7.769900959e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.37 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-6.020959369e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 3.139522843e-07 wvth0 = 2.037383109e-07 pvth0 = -1.921871807e-13
+ k1 = 0.64774
+ k2 = -1.159876940e-01 lk2 = 1.192792735e-07 wk2 = 6.507109893e-08 pk2 = -6.038447809e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 4.800372537e+04 lvsat = 1.113727084e-01 wvsat = 7.803562942e-02 pvsat = -1.147236904e-7
+ ua = -1.853319660e-09 lua = -1.149836434e-15 wua = -1.064060653e-15 pua = 1.184432712e-21
+ ub = 1.907761330e-18 lub = 1.237351967e-24 wub = 1.086473647e-24 pub = -1.274581413e-30
+ uc = 1.233672602e-10 luc = -6.760391057e-17 wuc = -6.054987076e-17 puc = 6.963797703e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 5.469807655e-03 lu0 = -2.995203876e-09 wu0 = -2.748005390e-09 pu0 = 2.951579426e-15
+ a0 = 4.389807499e-01 la0 = 1.132630777e-06 wa0 = 1.142815597e-06 pa0 = -1.270755774e-12
+ keta = -1.069159577e-02 lketa = -2.776228038e-09 wketa = -1.945222537e-09 pketa = 2.859759187e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.540930481e-01 lags = -5.229854616e-07 wags = -3.641351616e-07 pags = 5.530395492e-13
+ b0 = 2.309476920e-07 lb0 = -4.457151380e-13 wb0 = -2.378964461e-13 pb0 = 4.591258150e-19
+ b1 = 2.515816662e-07 lb1 = -7.412712717e-13 wb1 = -2.591512554e-13 pb1 = 7.635746418e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 6.079048215e-03 lpdiblc2 = 8.312278366e-09 wpdiblc2 = -1.403452963e-08 ppdiblc2 = 1.673432595e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -6.036893754e-02 ldelta = 1.231769098e-07 wdelta = 4.159331998e-08 pdelta = -6.017993903e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -2.415920654e-01 lkt1 = -4.133354721e-07 wkt1 = -3.084759394e-07 pkt1 = 3.496102953e-13
+ kt2 = -2.163859830e-01 lkt2 = 2.371946395e-07 wkt2 = 1.276890450e-07 pkt2 = -1.877214110e-13
+ at = 2.826925913e+05 lat = -4.749405954e-02 wat = 1.074051732e-01 pat = -1.734794315e-7
+ ute = -2.199431537e-01 lute = -1.432852348e-08 wute = 7.683332115e-08 pute = 1.272687532e-15
+ ua1 = 1.006505318e-09 lua1 = -4.563555278e-16 wua1 = -2.105477957e-16 pua1 = 3.095357891e-22
+ ub1 = -5.447551877e-19 lub1 = 6.216878428e-25 wub1 = 2.138662680e-25 pub1 = -3.144144246e-31
+ uc1 = 8.998935956e-11 luc1 = -1.469415214e-16 wuc1 = -1.029576660e-16 puc1 = 1.513626978e-22
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.38 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-3.746309694e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 9.327828330e-08 wvth0 = 5.924238548e-08 pvth0 = -5.200518110e-14
+ k1 = 0.64774
+ k2 = 1.072601287e-02 lk2 = -3.651395603e-09 wk2 = 4.025755349e-09 pk2 = -1.161643241e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.935178043e+05 lvsat = -2.979704770e-02 wvsat = -4.777871092e-02 pvsat = 7.334462801e-9
+ ua = -3.119231522e-09 lua = 7.828163018e-17 wua = 2.786832239e-16 pua = -1.182235457e-22
+ ub = 3.360330028e-18 lub = -1.718502928e-25 wub = -4.872864532e-25 pub = 2.521940801e-31
+ uc = 6.380530407e-11 luc = -9.820176640e-18 wuc = 8.310691709e-18 puc = 2.833246654e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.553981509e-03 lu0 = -1.664297195e-10 wu0 = 2.607962143e-10 pu0 = 3.260559361e-17
+ a0 = 2.023736329e+00 la0 = -4.048119250e-07 wa0 = -3.241178744e-07 pa0 = 1.523823981e-13
+ keta = -1.355325876e-02 wketa = 1.002542165e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 2.761343539e-01 lags = -1.563107242e-07 wags = 9.609560656e-08 pags = 1.065489706e-13
+ b0 = -7.062711487e-07 lb0 = 4.635230343e-13 wb0 = 5.678798412e-13 pb0 = -3.225940212e-19
+ b1 = -1.292305450e-06 lb1 = 7.565230944e-13 wb1 = 1.011198084e-12 pb1 = -4.688484181e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 1.521823935e-02 lpdiblc2 = -5.540622163e-10 wpdiblc2 = -2.815213474e-08 ppdiblc2 = 3.043044996e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 3.793411468e-02 ldelta = 2.780869525e-08 wdelta = -5.513016997e-09 pdelta = -1.447996174e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.636372778e-01 lkt1 = -3.890419475e-09 wkt1 = 6.811227264e-08 pkt1 = -1.573487560e-14
+ kt2 = 6.081379188e-02 lkt2 = -3.172933614e-08 wkt2 = -8.478148073e-08 pkt2 = 1.840580714e-14
+ at = 4.443537755e+05 lat = -2.043288491e-01 wat = -1.879219221e-01 pat = 1.130306734e-7
+ ute = -7.179722042e-02 lute = -1.580515599e-07 wute = -1.636009400e-08 pute = 9.168381328e-14
+ ua1 = -1.254155961e-11 lua1 = 5.322677053e-16 wua1 = 4.267774472e-16 pua1 = -3.087621087e-22
+ ub1 = 1.215403489e-18 lub1 = -1.085921297e-24 wub1 = -6.586241163e-25 pub1 = 5.320277593e-31
+ uc1 = -8.952938791e-11 luc1 = 2.721769391e-17 wuc1 = 6.933756358e-17 puc1 = -1.578865763e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.39 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 5.5e-07 wmax = 1.0e-6
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.010269380e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -3.535528401e-08 wvth0 = -7.669843389e-08 pvth0 = 1.190671542e-14
+ k1 = 0.64774
+ k2 = -5.946480726e-02 lk2 = 2.934846753e-08 wk2 = 2.473199205e-08 pk2 = -1.089657690e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.760051638e+05 lvsat = -2.156356735e-02 wvsat = -5.827588104e-02 pvsat = 1.226965484e-8
+ ua = -3.086907407e-09 lua = 6.308460889e-17 wua = 2.533804353e-16 pua = -1.063275662e-22
+ ub = 2.646268170e-18 lub = 1.638623191e-25 wub = -8.123619081e-26 pub = 6.129157951e-32
+ uc = 1.477477987e-11 luc = 1.323127916e-17 wuc = 4.332675812e-17 puc = -1.362938189e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.335555779e-03 lu0 = 4.064070455e-10 wu0 = 7.017805233e-10 pu0 = -1.747209744e-16
+ a0 = 1.1627
+ keta = -1.724188142e-02 lketa = 1.734187501e-09 wketa = 3.142267908e-09 pketa = -1.005981359e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -7.745090768e-01 lags = 3.376440316e-07 wags = 1.062503918e-06 pags = -3.478030652e-13
+ b0 = 9.047149019e-07 lb0 = -2.938740025e-13 wb0 = -3.870951670e-13 pb0 = 1.263827040e-19
+ b1 = -5.503158191e-09 lb1 = 1.515394310e-13 wb1 = 6.229700437e-13 pb1 = -2.863249461e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = 0.030097
+ pdiblc1 = 0.0
+ pdiblc2 = 2.042206481e-03 lpdiblc2 = 5.640583756e-09 wpdiblc2 = -4.474454554e-08 ppdiblc2 = 3.823128893e-14
+ pdiblcb = -0.025
+ drout = 0.43496
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.523937529e-01 ldelta = -2.600393139e-08 wdelta = -7.153664808e-08 pdelta = 1.656071830e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.940860710e-01 lkt1 = 5.743942839e-08 wkt1 = 1.369258638e-07 pkt1 = -4.808724140e-14
+ kt2 = 1.612187880e-01 lkt2 = -7.893424303e-08 wkt2 = -1.430252141e-07 pkt2 = 4.578880717e-14
+ at = -5.542513391e+04 lat = 3.063970628e-02 wat = 2.013034159e-01 pat = -6.996167316e-8
+ ute = -8.254924889e-01 lute = 1.962945021e-07 wute = 5.599479792e-07 pute = -1.792645458e-13
+ ua1 = 1.965680628e-09 lua1 = -3.977835649e-16 wua1 = -7.207655050e-16 pua1 = 2.307494726e-22
+ ub1 = -2.933875434e-18 lub1 = 8.648414428e-25 wub1 = 1.482526161e-24 pub1 = -4.746233378e-31
+ uc1 = -1.631896678e-10 luc1 = 6.184870619e-17 wuc1 = 1.120670080e-16 puc1 = -3.587769228e-23
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.40 pmos
* DC IV MOS Parameters
+ lmin = 2.0e-05 lmax = 1.0e-04 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.840824378e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} wvth0 = -6.853830342e-8
+ k1 = 0.64774
+ k2 = 2.963619883e-02 wk2 = -1.861977996e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.390670400e-09 wua = 2.088725182e-16
+ ub = 3.746938677e-18 wub = -3.886233872e-25
+ uc = 5.985726708e-11 wuc = 1.205033759e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.780762388e-03 wu0 = 2.393980317e-10
+ a0 = 2.077392191e+00 wa0 = -2.050565780e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.530359440e-01 wags = -2.253212290e-7
+ b0 = 4.767322002e-07 wb0 = -2.427420004e-13
+ b1 = 2.244393169e-07 wb1 = -4.820135035e-15
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.471549993e-03 wpdiblc2 = -6.024967955e-10
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.952522708e-03 wdelta = 2.100775520e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.822829231e-01 wkt1 = 1.205033759e-7
+ kt2 = -0.055045
+ at = 2.546853877e+05 wat = 1.596669730e-2
+ ute = -6.620897015e-01 wute = 2.182115298e-7
+ ua1 = 6.8217e-10
+ ub1 = -6.177426338e-20 wub1 = -5.125410254e-26
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.41 pmos
* DC IV MOS Parameters
+ lmin = 8e-06 lmax = 2.0e-05 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-6.913353782e-02+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -2.295546200e-06 wvth0 = -1.352187809e-07 pvth0 = 1.331618804e-12
+ k1 = 0.64774
+ k2 = 6.601476163e-02 lk2 = -7.264851741e-07 wk2 = -3.972254770e-08 pk2 = 4.214253316e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.390670400e-09 wua = 2.088725182e-16
+ ub = 3.746938677e-18 wub = -3.886233872e-25
+ uc = 5.985726708e-11 wuc = 1.205033759e-19
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.721517300e-03 lu0 = 1.183132998e-09 wu0 = 2.737653963e-10 pu0 = -6.863212544e-16
+ a0 = 1.689001593e+00 la0 = 7.756216555e-06 wa0 = 2.024414714e-08 pa0 = -4.499288149e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 6.530359440e-01 wags = -2.253212290e-7
+ b0 = 7.567643508e-07 lb0 = -5.592282650e-12 wb0 = -4.051852905e-13 pb0 = 3.244016058e-18
+ b1 = 2.552990080e-07 lb1 = -6.162725054e-13 wb1 = -2.272147151e-14 pb1 = 3.574922851e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 3.978198536e-03 lpdiblc2 = -5.005813487e-08 wpdiblc2 = -2.056573536e-09 ppdiblc2 = 2.903812334e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.278619900e-02 ldelta = -2.562903765e-07 wdelta = -5.343886096e-09 pdelta = 1.486709719e-13
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -8.822829231e-01 wkt1 = 1.205033759e-7
+ kt2 = -0.055045
+ at = 2.169271070e+05 lat = 7.540383412e-01 wat = 3.786982286e-02 pat = -4.374085933e-7
+ ute = -6.620897015e-01 wute = 2.182115298e-7
+ ua1 = 6.8217e-10
+ ub1 = -3.090260684e-21 lub1 = -1.171928043e-24 wub1 = -8.529598830e-26 pub1 = 6.798213947e-31
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.42 pmos
* DC IV MOS Parameters
+ lmin = 4e-06 lmax = 8e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-5.354722059e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 1.421240604e-06 wvth0 = 1.184842370e-07 pvth0 = -6.904310358e-13
+ k1 = 0.64774
+ k2 = -9.021295151e-02 lk2 = 5.186723527e-07 wk2 = 4.363202153e-08 pk2 = -2.429226715e-13
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.452731505e-09 lua = 4.946360063e-16 wua = 2.680764828e-16 pua = -4.718641821e-22
+ ub = 4.131138935e-18 lub = -3.062131769e-24 wub = -6.292267045e-25 pub = 1.917643326e-30
+ uc = 1.044628759e-10 luc = -3.555131700e-16 wuc = -2.264212529e-17 puc = 1.814214510e-22
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 2.470849677e-03 lu0 = -4.789154698e-09 wu0 = -1.190027203e-10 pu0 = 2.444097587e-15
+ a0 = 3.047256683e+00 la0 = -3.069273462e-06 wa0 = -7.477996680e-07 pa0 = 1.622132424e-12
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.702249165e-01 lags = -9.340131031e-07 wags = -2.780665792e-07 pags = 4.203880895e-13
+ b0 = -4.100456838e-07 lb0 = 3.707362513e-12 wb0 = 2.484670254e-13 pb0 = -1.965687679e-18
+ b1 = 2.506781471e-07 lb1 = -5.794435742e-13 wb1 = -9.602466354e-15 pb1 = 2.529319118e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 1.956862042e-03 lpdiblc2 = -3.394778992e-08 wpdiblc2 = -2.406429253e-09 ppdiblc2 = 3.182652414e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -5.606173076e-03 ldelta = -2.999905415e-08 wdelta = 8.547366508e-09 pdelta = 3.795567445e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.015130388e+00 lkt1 = 1.058813559e-06 wkt1 = 1.803053603e-07 pkt1 = -4.766304870e-13
+ kt2 = -0.055045
+ at = 3.534943989e+05 lat = -3.344227774e-01 wat = -3.389515349e-02 pat = 1.345686742e-7
+ ute = -1.224206355e+00 lute = 4.480151237e-06 wute = 4.347943833e-07 pute = -1.726196747e-12
+ ua1 = 6.683538954e-10 lua1 = 1.101163570e-16
+ ub1 = -1.781691491e-19 lub1 = 2.234760837e-25
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.43 pmos
* DC IV MOS Parameters
+ lmin = 2e-06 lmax = 4e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.848812235e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = 2.934356816e-08 wvth0 = -5.704776345e-08 pvth0 = 6.456458215e-15
+ k1 = 0.64774
+ k2 = 4.630594560e-02 lk2 = -2.332746405e-08 wk2 = -1.887691093e-08 pk2 = 5.246854121e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.284186546e-09 lua = -1.745119185e-16 wua = 1.294392535e-16 pua = 7.854572038e-23
+ ub = 3.271937167e-18 lub = 3.490238370e-25 wub = -1.066425755e-25 pub = -1.570914408e-31
+ uc = 1.491622960e-11 wuc = 2.305430420e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.484154372e-03 lu0 = -8.718312660e-10 wu0 = 3.489104397e-10 pu0 = 5.864144938e-16
+ a0 = 2.043616137e+00 la0 = 9.153250365e-07 wa0 = -2.054765302e-07 pa0 = -5.309690697e-13
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 3.661894890e-01 lags = 6.700661291e-07 wags = -1.205427559e-07 pags = -2.050043302e-13
+ b0 = 8.321360521e-07 lb0 = -1.224279095e-12 wb0 = -4.012254284e-13 pb0 = 6.136855679e-19
+ b1 = 1.390496184e-07 lb1 = -1.362621290e-13 wb1 = 3.535069502e-14 pb1 = 7.446134292e-20
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -1.854234674e-02 lpdiblc2 = 4.743704132e-08 wpdiblc2 = 1.020706666e-08 ppdiblc2 = -1.825088359e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = -5.465529581e-02 ldelta = 1.647330752e-07 wdelta = 3.846349454e-08 pdelta = -8.081569170e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -6.987449933e-01 lkt1 = -1.972823340e-07 wkt1 = 3.142626353e-08 pkt1 = 1.144411146e-13
+ kt2 = -0.055045
+ at = 3.058455927e+05 lat = -1.452501077e-1
+ ute = -1.480090102e-01 lute = 2.074917287e-07 wute = 3.031714507e-08 pute = -1.203634619e-13
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.44 pmos
* DC IV MOS Parameters
+ lmin = 1.5e-06 lmax = 2e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.699871075e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} wvth0 = -5.377061471e-8
+ k1 = 0.64774
+ k2 = 3.446546480e-02 wk2 = -1.621372922e-8
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 123760.0
+ ua = -3.372764757e-09 wua = 1.693072431e-16
+ ub = 3.449093588e-18 wub = -1.863785547e-25
+ uc = 1.491622960e-11 wuc = 2.305430420e-17
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.041633001e-03 wu0 = 6.465608633e-10
+ a0 = 2.508213938e+00 wa0 = -4.749841399e-7
+ keta = -0.01258
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 7.062995465e-01 wags = -2.245982087e-7
+ b0 = 2.107203212e-07 wb0 = -8.973283885e-14
+ b1 = 6.988611569e-08 wb1 = 7.314554916e-14
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = 5.535597434e-03 wpdiblc2 = 9.433405942e-10
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.895940018e-02 wdelta = -2.556679958e-9
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -7.988809397e-01 wkt1 = 8.951392438e-8
+ kt2 = -0.055045
+ at = 232120.0
+ ute = -4.269101145e-02 wute = -3.077656220e-8
+ ua1 = 6.9609e-10
+ ub1 = -1.2188e-19
+ uc1 = -9.961e-12
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 3.0e-6
+ sbref = 3.0e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.45 pmos
* DC IV MOS Parameters
+ lmin = 1e-06 lmax = 1.5e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.362415621e-02+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -2.298762110e-07 wvth0 = -1.376271075e-07 pvth0 = 1.232812035e-13
+ k1 = 0.64774
+ k2 = 8.157365228e-02 lk2 = -6.925586628e-08 wk2 = -4.953186729e-08 pk2 = 4.898249408e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 3.859932583e+05 lvsat = -3.855209136e-01 wvsat = -1.180280428e-01 pvsat = 1.735183369e-7
+ ua = -4.552513411e-09 lua = 1.734401585e-15 wua = 5.017092521e-16 pua = -4.886791515e-22
+ ub = 5.301110960e-18 lub = -2.722734080e-24 wub = -8.819677529e-25 pub = 1.022616982e-30
+ uc = -8.626031317e-11 luc = 1.487441885e-16 wuc = 6.105256902e-17 puc = -5.586295904e-23
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = -1.887923944e-04 lu0 = 1.808903743e-09 wu0 = 5.344805953e-10 pu0 = 1.647742456e-16
+ a0 = 4.615072939e+00 la0 = -3.097388226e-06 wa0 = -1.279685369e-06 pa0 = 1.183027489e-12
+ keta = -1.911678388e-02 lketa = 9.610020131e-09 wketa = 2.942127981e-09 pketa = -4.325354741e-15
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = -9.686185723e-01 lags = 2.462372498e-06 wags = 5.771803768e-07 pags = -1.178730779e-12
+ b0 = -7.407497322e-07 lb0 = 1.398798942e-12 wb0 = 3.257735693e-13 pb0 = -6.108546683e-19
+ b1 = -6.202082953e-08 lb1 = 1.939223360e-13 wb1 = -7.723421083e-14 pb1 = 2.210800522e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -5.061066833e-01 wpclm = 3.110453222e-7
+ pdiblc1 = 0.0
+ pdiblc2 = -4.650897517e-02 lpdiblc2 = 7.651306819e-08 wpdiblc2 = 1.647115168e-08 ppdiblc2 = -2.282813382e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 2.050977276e-02 ldelta = 1.242217752e-08 wdelta = -5.323449318e-09 pdelta = 4.067552140e-15
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -1.205857425e+00 lkt1 = 5.983144451e-07 wkt1 = 2.508828246e-07 pkt1 = -2.372356819e-13
+ kt2 = 3.734145260e-03 lkt2 = -8.641386651e-8
+ at = 1.013121694e+06 lat = -1.148185736e+00 wat = -3.163079844e-01 pat = 4.650186017e-7
+ ute = -1.867676258e-01 lute = 2.118135142e-07 wute = 5.758859555e-08 pute = -1.299095948e-13
+ ua1 = 3.520658619e-10 lua1 = 5.057653666e-16 wua1 = 1.690846796e-16 pua1 = -2.485789963e-22
+ ub1 = -4.789907938e-19 lub1 = 5.250046480e-25 wub1 = 1.757171324e-25 pub1 = -2.583296635e-31
+ uc1 = -8.749692869e-11 luc1 = 1.139890579e-16 puc1 = 1.175494351e-38
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 2.74e-6
+ sbref = 2.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.46 pmos
* DC IV MOS Parameters
+ lmin = 5e-07 lmax = 1e-06 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope2/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.804498169e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope2/sqrt(1))} lvth0 = -6.803113043e-08 wvth0 = -5.339977088e-08 pvth0 = 4.156847409e-14
+ k1 = 0.64774
+ k2 = 3.001954362e-02 lk2 = -1.924090554e-08 wk2 = -7.166190316e-09 pk2 = 7.881644398e-15
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = 1.493031557e+05 lvsat = -1.558971940e-01 wvsat = -2.213032387e-02 pvsat = 8.048364444e-8
+ ua = -2.773386508e-09 lua = 8.390516121e-18 wua = 7.806268138e-17 pua = -7.768054915e-23
+ ub = 2.101841368e-18 lub = 3.810213183e-25 wub = 2.427477163e-25 pub = -6.852010704e-32
+ uc = 8.818247204e-11 luc = -2.049060739e-17 wuc = -5.830210901e-18 puc = 9.023035485e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 8.976596231e-04 lu0 = 7.548877507e-10 wu0 = 1.221608664e-09 pu0 = -5.018396151e-16
+ a0 = 3.381192980e+00 la0 = -1.900345753e-06 wa0 = -1.111562188e-06 pa0 = 1.019923625e-12
+ keta = -9.211027385e-03 wketa = -1.516334147e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 1.443657067e+00 lags = 1.221153479e-07 wags = -5.811703089e-07 pags = -5.496265270e-14
+ b0 = 1.097637196e-06 lb0 = -3.847029446e-13 wb0 = -4.785457425e-13 pb0 = 1.694516904e-19
+ b1 = -4.770794506e-07 lb1 = 5.965893819e-13 wb1 = 5.382952646e-13 pb1 = -3.760727907e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -9.035364757e-01 lpclm = 3.855645260e-07 wpclm = 5.415895756e-07 ppclm = -2.236613547e-13
+ pdiblc1 = 0.0
+ pdiblc2 = -1.269624624e-01 lpdiblc2 = 1.545646166e-07 wpdiblc2 = 5.432518420e-08 ppdiblc2 = -5.955203420e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 9.822717640e-02 ldelta = -6.297497304e-08 wdelta = -4.048829859e-08 pdelta = 3.818255483e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -4.571521952e-01 lkt1 = -1.280381901e-07 wkt1 = -5.166724596e-08 pkt1 = 5.628175637e-14
+ kt2 = -0.085339
+ at = -3.394197285e+05 lat = 1.639755627e-01 wat = 2.667356822e-01 pat = -1.006182962e-7
+ ute = 1.552726718e-01 lute = -1.200151703e-07 wute = -1.480806136e-07 pute = 6.961936009e-14
+ ua1 = 9.204698604e-10 lua1 = -4.566893058e-17 wua1 = -1.144512814e-16 pua1 = 2.649199860e-23
+ ub1 = 9.346713997e-19 lub1 = -8.464526608e-25 wub1 = -4.957748000e-25 pub1 = 3.931148772e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.74e-6
+ sbref = 1.74e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.model sky130_fd_pr__pfet_01v8_lvt.47 pmos
* DC IV MOS Parameters
+ lmin = 3.5e-07 lmax = 5e-07 wmin = 4.2e-07 wmax = 5.5e-7
+ level = 54.0
+ tnom = 30.0
+ version = 4.5
+ toxm = 4.23e-9
+ xj = 1.5e-7
+ lln = 1.0
+ lwn = 1.0
+ wln = 1.0
+ wwn = 1.0
+ lint = 1.49275e-8
+ ll = 0.0
+ lw = 0.0
+ lwl = 0.0
+ wint = -1.5044e-8
+ wl = 0.0
+ ww = 0.0
+ wwl = 0.0
+ xl = 0.0
+ xw = 0.0
+ mobmod = 0.0
+ binunit = 2.0
+ dwg = -7.916e-9
+ dwb = 0.0
* BSIM4 - Model Selectors
+ igcmod = 0.0
+ igbmod = 0.0
+ rgatemod = 0.0
+ rbodymod = 1.0
+ trnqsmod = 0.0
+ acnqsmod = 0.0
+ fnoimod = 1.0
+ tnoimod = 1.0
+ permod = 1.0
+ geomod = 0.0
+ rdsmod = 0.0
+ tempmod = 0.0
+ lintnoi = 0.0
+ vfbsdoff = 0.0
+ lambda = 0.0
+ vtl = 0.0
+ lc = 5.0e-9
+ xn = 3.0
+ rnoia = 0.69
+ rnoib = 0.34
+ tnoia = 25000000.0
+ tnoib = 0.0
* BSIM4 - Process Parameters
+ epsrox = 3.9
+ toxe = {4.075605e-09+MC_MM_SWITCH*(4.075605e-09*(sky130_fd_pr__pfet_01v8_lvt__toxe_slope3/sqrt(1)))}
+ dtox = 0.0
+ ndep = 1.7000000000000000e+17
+ nsd = 1.0e+20
+ rshg = 0.1
+ rsh = 1.0
* Threshold Voltage Parameters
+ vth0 = {-1.097473764e-01+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__vth0_slope1/sqrt(1))} lvth0 = -1.012715293e-07 wvth0 = -7.163981225e-08 pvth0 = 5.014393834e-14
+ k1 = 0.64774
+ k2 = 3.139230846e-02 lk2 = -1.988630406e-08 wk2 = -2.797313049e-08 pk2 = 1.766392329e-14
+ k3 = 3.39
+ dvt0 = 2.4422
+ dvt1 = 0.16136
+ dvt2 = 0.026237
+ dvt0w = 0.5
+ dvt1w = 1928100.0
+ dvt2w = -0.032
+ w0 = 1.0e-8
+ k3b = 1.0
* NEW BSIM4 Parameters for Level 54
+ phin = 0.0
+ lpe0 = 0.0
+ lpeb = 0.0
+ vbm = -3.0
+ dvtp0 = 0.0
+ dvtp1 = 0.0
* Mobility Parameters
+ vsat = -5.712960980e+05 lvsat = 1.828889422e-01 wvsat = 3.752246133e-01 pvsat = -1.063307925e-7
+ ua = -2.063875741e-09 lua = -3.251824237e-16 wua = -3.400679578e-16 pua = 1.189014802e-22
+ ub = 1.314830304e-18 lub = 7.510306350e-25 wub = 6.911149380e-25 pub = -2.793177145e-31
+ uc = 7.614770502e-11 luc = -1.483252185e-17 wuc = 7.725060712e-18 puc = 2.650092313e-24
+ rdsw = 484.7
+ prwb = 0.1
+ prwg = 0.052
+ wr = 1.0
+ u0 = 1.718685900e-03 lu0 = 3.688863518e-10 wu0 = 4.795313376e-10 pu0 = -1.529556702e-16
+ a0 = -6.608488431e-01 wa0 = 1.057818801e-6
+ keta = -9.211027385e-03 wketa = -1.516334147e-9
+ a1 = 0.0
+ a2 = 0.46703705
+ ags = 4.189369878e+00 lags = -1.168767802e-06 wags = -1.816982697e-06 pags = 5.260483623e-13
+ b0 = 8.756379653e-07 lb0 = -2.803311164e-13 wb0 = -3.702279849e-13 pb0 = 1.185266382e-19
+ b1 = 2.481952424e-06 lb1 = -7.945846588e-13 wb1 = -8.199730901e-13 pb1 = 2.625102849e-19
* BSIM4 - Mobility Parameters
+ eu = 1.67
+ rdswmin = 0.0
+ rdw = 0.0
+ rdwmin = 0.0
+ rsw = 0.0
+ rswmin = 0.0
* Subthreshold Current Parameters
+ voff = {-0.1819+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__voff_slope/sqrt(1))}
+ nfactor = {2.5373+MC_MM_SWITCH*(sky130_fd_pr__pfet_01v8_lvt__nfactor_slope/sqrt(1))}
+ up = 0.0
+ ud = 0.0
+ lp = 1.0
+ tvfbsdoff = 0.0
+ tvoff = 0.0
+ cit = -6.393105e-11
+ cdsc = 2.8125e-7
+ cdscb = 1.0e-4
+ cdscd = 1.0e-10
+ eta0 = 0.2
+ etab = -0.00025
+ dsub = 1.0
* BSIM4 - Sub-threshold parameters
+ voffl = 0.0
+ minv = 0.0
* Rout Parameters
+ pclm = -8.343942911e-02 wpclm = 6.586112009e-8
+ pdiblc1 = 0.0
+ pdiblc2 = -5.498729596e-02 lpdiblc2 = 1.207258520e-07 wpdiblc2 = -1.166241553e-08 ppdiblc2 = -2.852829413e-14
+ pdiblcb = -0.025
+ drout = 4.650812738e-01 wdrout = -1.747298950e-8
+ pscbe1 = 800000000.0
+ pscbe2 = 8.6797e-9
+ pvag = 0.0
+ delta = 1.262736113e-01 ldelta = -7.616086416e-08 wdelta = -5.638466733e-08 pdelta = 4.565615312e-14
+ alpha0 = 5.0449517e-13
+ alpha1 = -4.0583656e-18
+ beta0 = 6.2016506
* BSIM4 - Rout Parameters
+ fprout = 0.0
+ pdits = 0.0
+ pditsl = 0.0
+ pditsd = 0.0
* BSIM4 - Gate Induced Drain Leakage Model Parameters
+ agidl = 0.0
+ bgidl = 2300000000.0
+ cgidl = 0.5
+ egidl = 0.8
* BSIM4 - Gate Leakage Current Parameters
+ aigbacc = 0.43
+ bigbacc = 0.054
+ cigbacc = 0.075
+ nigbacc = 1.0
+ aigbinv = 0.35
+ bigbinv = 0.03
+ cigbinv = 0.006
+ eigbinv = 1.1
+ nigbinv = 3.0
+ aigc = 0.43
+ bigc = 0.054
+ cigc = 0.075
+ nigc = 1.0
+ aigsd = 0.43
+ bigsd = 0.054
+ cigsd = 0.075
+ dlcig = 0.0
+ poxedge = 1.0
+ pigcd = 1.0
+ ntox = 1.0
+ toxref = 4.23e-9
* Temperature Effects Parameters
+ kt1 = -9.256957515e-01 lkt1 = 9.224522017e-08 wkt1 = 2.132710601e-07 pkt1 = -6.827766354e-14
+ kt2 = -0.085339
+ at = 6.742000300e+03 lat = 1.229356704e-03 wat = 1.652410073e-01 pat = -5.290108229e-8
+ ute = 1.397886050e-01 lute = -1.127354137e-7
+ ua1 = 1.037107415e-09 lua1 = -1.005054938e-16 wua1 = -1.821113273e-16 pua1 = 5.830203088e-23
+ ub1 = -2.217316449e-18 lub1 = 6.354386665e-25 wub1 = 1.066858892e-24 pub1 = -3.415495401e-31
+ uc1 = 3.0e-11
+ kt1l = 0.0
+ prt = 0.0
* BSIM4 - High Speed RF Model Parameters
+ xrcrg1 = 12.0
+ xrcrg2 = 1.0
+ rbpb = 50.0
+ rbpd = 50.0
+ rbps = 50.0
+ rbdb = 50.0
+ rbsb = 50.0
+ gbmin = 1.0e-12
* BSIM4 - Flicker and Thermal Noise Parameters
+ noia = 3.0e+41
+ noib = 0.0
+ noic = 0.0
+ em = 41000000.0
+ af = 1.0
+ ef = 0.88
+ kf = 0.0
+ ntnoi = 1.0
* BSIM4 - Layout Dependent Parasitic Model Parameters
+ dmcg = 0.0
+ dmcgt = 0.0
+ dmdg = 0.0
+ xgw = 0.0
+ xgl = 0.0
+ ngcon = 1.0
* Diode DC IV Parameters
* BSIM4 - Diode DC IV parameters
+ diomod = 1.0
+ njs = 1.3632
+ jss = 2.1483e-5
+ jsws = 1.4472e-10
+ xtis = 5.2
+ bvs = 12.69
+ xjbvs = 1.0
+ ijthsrev = 0.1
+ ijthsfwd = 0.1
* Diode and FET Capacitance Parameters
+ tpb = 0.001671
+ tpbsw = 0.001246
+ tpbswg = 0.0
+ tcj = 0.0012407
+ tcjsw = 0.00037357
+ tcjswg = 2.0e-12
+ cgdo = 7.24e-11
+ cgso = 7.24e-11
+ cgbo = 1.0e-13
+ capmod = 2.0
+ xpart = 0.0
+ cgsl = 0.0
+ cgdl = 0.0
+ cf = 0.0
+ clc = 7.0e-8
+ cle = 0.492
+ dlc = 2.0382e-8
+ dwc = -2.252e-8
+ vfbcv = -1.0
+ acde = 0.44
+ moin = 8.7
+ noff = 2.6123
+ voffcv = 0.112
+ ngate = 1.0e+23
+ lwc = 0.0
+ llc = 0.0
+ lwlc = 0.0
+ wlc = 0.0
+ wwc = 0.0
+ wwlc = 0.0
* BSIM4 - FET and Diode capacitance parameters
+ ckappas = 0.6
+ cjs = 0.0007144615823
+ mjs = 0.3362
+ pbs = 0.6587
+ cjsws = 8.55153728e-11
+ mjsws = 0.2659
+ pbsws = 0.7418
+ cjswgs = 2.232631466e-10
+ mjswgs = 0.9274
+ pbswgs = 1.4338
* Stress Parameters
+ saref = 1.44e-6
+ sbref = 1.44e-6
+ wlod = {0+sky130_fd_pr__pfet_01v8_lvt__wlod_diff}
+ kvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__kvth0_diff}
+ lkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__lkvth0_diff}
+ wkvth0 = {0+sky130_fd_pr__pfet_01v8_lvt__wkvth0_diff}
+ pkvth0 = 0.0
+ llodvth = 0.0
+ wlodvth = 1.0
+ stk2 = 0.0
+ lodk2 = 1.0
+ lodeta0 = 1.0
+ ku0 = {0+sky130_fd_pr__pfet_01v8_lvt__ku0_diff}
+ lku0 = {0+sky130_fd_pr__pfet_01v8_lvt__lku0_diff}
+ wku0 = {0+sky130_fd_pr__pfet_01v8_lvt__wku0_diff}
+ pku0 = 0.0
+ llodku0 = 0.0
+ wlodku0 = 1.0
+ kvsat = {0+sky130_fd_pr__pfet_01v8_lvt__kvsat_diff}
+ steta0 = 0.0
+ tku0 = 0.0
.ends sky130_fd_pr__pfet_01v8_lvt
