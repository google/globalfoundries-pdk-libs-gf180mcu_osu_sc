magic
tech gf180mcuC
timestamp 1659392489
<< nwell >>
rect 0 97 44 159
<< metal1 >>
rect 0 147 44 159
rect 0 -3 44 9
<< end >>
