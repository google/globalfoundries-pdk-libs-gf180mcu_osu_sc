# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__tinv_2
  CLASS CORE ;
  ORIGIN 3.3 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__tinv_2 -3.3 0 ;
  SIZE 6.5 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT -3.3 5.55 3.2 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
        RECT -2.2 3.5 -1.95 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT -3.3 0 3.2 0.6 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
        RECT -2.2 0 -1.95 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -1.35 1.45 -1.05 2.9 ;
      LAYER MET2 ;
        RECT -1.45 1.5 -0.95 1.9 ;
      LAYER VIA12 ;
        RECT -1.33 1.57 -1.07 1.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -2.85 2.2 -2.35 2.5 ;
      LAYER MET2 ;
        RECT -2.85 2.15 -2.35 2.55 ;
      LAYER VIA12 ;
        RECT -2.73 2.22 -2.47 2.48 ;
    END
  END EN
  PIN EN_BAR
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT -2.15 2.85 -1.65 3.15 ;
      LAYER MET2 ;
        RECT -2.15 2.8 -1.65 3.2 ;
      LAYER VIA12 ;
        RECT -2.03 2.87 -1.77 3.13 ;
    END
  END EN_BAR
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.4 3 2.65 3.25 ;
        RECT 2.4 2.05 2.65 3.25 ;
        RECT 1.4 2.05 2.65 2.3 ;
        RECT 1.4 3 1.95 3.9 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 1.55 3.5 2.05 3.8 ;
        RECT 1.6 3.45 2 3.85 ;
      LAYER VIA12 ;
        RECT 1.67 3.52 1.93 3.78 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT -0.9 2.8 0.65 3.2 ;
    LAYER VIA12 ;
      RECT 0.27 2.87 0.53 3.13 ;
      RECT -0.78 2.87 -0.52 3.13 ;
    LAYER MET1 ;
      RECT -0.3 3.5 -0.05 5.2 ;
      RECT -0.25 2.2 0 3.7 ;
      RECT 0.85 2.1 1.1 2.55 ;
      RECT -0.3 0.95 -0.05 2.55 ;
      RECT -0.3 2.2 1.1 2.45 ;
      RECT -0.8 0.95 -0.55 5.2 ;
      RECT -0.8 2.75 -0.5 3.25 ;
      RECT 0.25 2.75 0.55 3.25 ;
  END
END gf180mcu_osu_sc_gp9t3v3__tinv_2
