magic
tech gf180mcuC
timestamp 1659394356
<< nwell >>
rect 0 97 88 159
<< metal1 >>
rect 0 147 88 159
rect 0 -3 88 9
<< end >>
