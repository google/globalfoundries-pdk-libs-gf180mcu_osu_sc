# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__inv_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__inv_4 0 0 ;
  SIZE 4.8 BY 6.15 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp9t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.8 6.15 ;
        RECT 4 3.5 4.25 6.15 ;
        RECT 2.25 3.5 2.5 6.15 ;
        RECT 0.55 3.5 0.8 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 3.95 0 4.2 1.8 ;
        RECT 2.25 0 2.5 1.8 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.4 2.2 0.9 2.5 ;
      LAYER MET2 ;
        RECT 0.4 2.15 0.9 2.55 ;
      LAYER VIA12 ;
        RECT 0.52 2.22 0.78 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 3.5 3.75 3.8 ;
        RECT 3.1 0.95 3.35 5.2 ;
        RECT 1.4 3 3.35 3.25 ;
        RECT 1.4 2.05 3.35 2.3 ;
        RECT 1.4 0.95 1.65 5.2 ;
      LAYER MET2 ;
        RECT 3.25 3.5 3.75 3.8 ;
        RECT 3.3 3.45 3.7 3.85 ;
      LAYER VIA12 ;
        RECT 3.37 3.52 3.63 3.78 ;
    END
  END Y
END gf180mcu_osu_sc_gp9t3v3__inv_4
