* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp12t3v3__dffsrn_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp12t3v3__dffsrn_1 D Q QN CLK RN SN VDD VSS
X0 a_156_109# a_133_14# a_82_14# VDD pmos_3p3 w=1.7u l=0.3u
X1 VSS a_41_109# a_156_19# VSS nmos_3p3 w=0.85u l=0.3u
X2 a_82_14# a_133_81# a_123_109# VDD pmos_3p3 w=1.7u l=0.3u
X3 a_212_109# a_133_81# a_195_19# VDD pmos_3p3 w=1.7u l=0.3u
X4 VDD CLK a_133_81# VDD pmos_3p3 w=1.7u l=0.3u
X5 a_195_19# a_133_81# a_184_19# VSS nmos_3p3 w=0.85u l=0.3u
X6 a_133_14# a_133_81# VSS VSS nmos_3p3 w=0.85u l=0.3u
X7 a_25_19# RN VDD VDD pmos_3p3 w=1.7u l=0.3u
X8 a_123_109# D VDD VDD pmos_3p3 w=1.7u l=0.3u
X9 a_41_109# a_25_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X10 VSS a_216_68# QN VSS nmos_3p3 w=0.85u l=0.3u
X11 Q QN VDD VDD pmos_3p3 w=1.7u l=0.3u
X12 a_310_19# a_195_19# VSS VSS nmos_3p3 w=0.85u l=0.3u
X13 VDD a_216_68# QN VDD pmos_3p3 w=1.7u l=0.3u
X14 a_25_19# RN VSS VSS nmos_3p3 w=0.85u l=0.3u
X15 a_82_14# a_133_14# a_123_19# VSS nmos_3p3 w=0.85u l=0.3u
X16 VSS CLK a_133_81# VSS nmos_3p3 w=0.85u l=0.3u
X17 a_216_68# SN a_310_19# VSS nmos_3p3 w=0.85u l=0.3u
X18 a_212_19# a_133_14# a_195_19# VSS nmos_3p3 w=0.85u l=0.3u
X19 VSS a_216_68# a_212_19# VSS nmos_3p3 w=0.85u l=0.3u
X20 a_77_19# SN a_41_109# VSS nmos_3p3 w=0.85u l=0.3u
X21 a_57_109# a_82_14# VDD VDD pmos_3p3 w=1.7u l=0.3u
X22 Q QN VSS VSS nmos_3p3 w=0.85u l=0.3u
X23 a_216_68# a_25_19# a_291_109# VDD pmos_3p3 w=1.7u l=0.3u
X24 a_57_109# a_25_19# a_41_109# VDD pmos_3p3 w=1.7u l=0.3u
X25 VDD SN a_57_109# VDD pmos_3p3 w=1.7u l=0.3u
X26 a_195_19# a_133_14# a_184_109# VDD pmos_3p3 w=1.7u l=0.3u
X27 a_291_109# SN VDD VDD pmos_3p3 w=1.7u l=0.3u
X28 VDD a_195_19# a_291_109# VDD pmos_3p3 w=1.7u l=0.3u
X29 a_184_109# a_41_109# VDD VDD pmos_3p3 w=1.7u l=0.3u
X30 VSS a_82_14# a_77_19# VSS nmos_3p3 w=0.85u l=0.3u
X31 a_156_19# a_133_81# a_82_14# VSS nmos_3p3 w=0.85u l=0.3u
X32 VDD a_41_109# a_156_109# VDD pmos_3p3 w=1.7u l=0.3u
X33 a_133_14# a_133_81# VDD VDD pmos_3p3 w=1.7u l=0.3u
X34 a_123_19# D VSS VSS nmos_3p3 w=0.85u l=0.3u
X35 VDD a_216_68# a_212_109# VDD pmos_3p3 w=1.7u l=0.3u
X36 a_184_19# a_41_109# VSS VSS nmos_3p3 w=0.85u l=0.3u
X37 VSS a_25_19# a_216_68# VSS nmos_3p3 w=0.85u l=0.3u
.ends
