magic
tech gf180mcuC
timestamp 1660766026
<< nwell >>
rect 0 97 32 159
<< metal1 >>
rect 0 147 32 159
rect 0 36 32 48
<< labels >>
rlabel metal1 10 153 10 153 1 VDD
rlabel metal1 6 42 6 42 1 GND
<< end >>
