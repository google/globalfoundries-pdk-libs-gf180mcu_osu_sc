* Copyright 2022 Google LLC
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*      http://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__aoi22_1.ext - technology: gf180mcuC

.subckt gf180mcu_osu_sc_gp9t3v3__aoi22_1 A0 A1 B0 B1 Y VDD VSS
X0 a_9_70# A1 VDD VDD pmos_3p3 w=1.7u l=0.3u
X1 a_56_19# B0 Y VSS nmos_3p3 w=0.85u l=0.3u
X2 Y B0 a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X3 VDD A0 a_9_70# VDD pmos_3p3 w=1.7u l=0.3u
X4 VSS B1 a_56_19# VSS nmos_3p3 w=0.85u l=0.3u
X5 a_28_19# A0 VSS VSS nmos_3p3 w=0.85u l=0.3u
X6 a_9_70# B1 Y VDD pmos_3p3 w=1.7u l=0.3u
X7 Y A1 a_28_19# VSS nmos_3p3 w=0.85u l=0.3u
.ends
