

.option scale=0.05u

.subckt gf180mcu_osu_sc_12T_fill_2
.ends

