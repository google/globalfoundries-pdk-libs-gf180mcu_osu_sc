# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp9t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__oai31_1 0 0 ;
  SIZE 4.9 BY 6.15 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 5.55 4.9 6.15 ;
        RECT 3.95 4.45 4.2 6.15 ;
        RECT 1 3.5 1.25 6.15 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.9 0.6 ;
        RECT 2.25 0 2.5 1.4 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.75 2.2 2.25 2.5 ;
      LAYER MET2 ;
        RECT 1.75 2.15 2.25 2.55 ;
      LAYER VIA12 ;
        RECT 1.87 2.22 2.13 2.48 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 2.85 3.05 3.15 ;
      LAYER MET2 ;
        RECT 2.55 2.8 3.05 3.2 ;
      LAYER VIA12 ;
        RECT 2.67 2.87 2.93 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.75 2.2 1.25 2.5 ;
      LAYER MET2 ;
        RECT 0.75 2.15 1.25 2.55 ;
      LAYER VIA12 ;
        RECT 0.87 2.22 1.13 2.48 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.25 2.2 3.75 2.5 ;
      LAYER MET2 ;
        RECT 3.25 2.15 3.75 2.55 ;
      LAYER VIA12 ;
        RECT 3.37 2.22 3.63 2.48 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 3.5 4.4 3.8 ;
        RECT 4 3.45 4.35 3.8 ;
        RECT 4.05 0.95 4.3 3.8 ;
        RECT 3 3.5 3.35 5.2 ;
      LAYER MET2 ;
        RECT 3.9 3.5 4.4 3.8 ;
        RECT 3.95 3.45 4.35 3.85 ;
      LAYER VIA12 ;
        RECT 4.02 3.52 4.28 3.78 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.65 3.45 1.9 ;
      RECT 3.1 0.95 3.45 1.9 ;
      RECT 1.4 0.95 1.65 1.9 ;
  END
END gf180mcu_osu_sc_gp9t3v3__oai31_1
