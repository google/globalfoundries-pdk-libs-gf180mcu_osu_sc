# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_lshifup
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_12T_lshifup 0 0 ;
  SIZE 6.6 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF180_3p3_12t ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 1.85 8.1 ;
        RECT 0.55 5.45 0.85 8.1 ;
    END
  END VDD
  PIN VDDH
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER MET1 ;
        RECT 2.1 7.5 6.6 8.1 ;
        RECT 4.85 5.45 5.15 8.1 ;
        RECT 3.15 5.45 3.45 8.1 ;
    END
  END VDDH
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 6.6 0.6 ;
        RECT 4.85 0 5.15 1.8 ;
        RECT 3.15 0 3.45 1.8 ;
        RECT 0.55 0 0.85 1.8 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.8 2.2 3.3 2.5 ;
        RECT 0.6 2.2 1.1 2.5 ;
      LAYER MET2 ;
        RECT 2.8 2.15 3.3 2.55 ;
        RECT 0.6 2.2 3.3 2.5 ;
        RECT 0.6 2.15 1.1 2.55 ;
      LAYER VIA12 ;
        RECT 0.72 2.22 0.98 2.48 ;
        RECT 2.92 2.22 3.18 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 5.7 4.15 6.1 4.45 ;
        RECT 5.75 0.95 6.05 7.15 ;
      LAYER MET2 ;
        RECT 5.65 4.1 6.15 4.5 ;
      LAYER VIA12 ;
        RECT 5.77 4.17 6.03 4.43 ;
    END
  END Y
  OBS
    LAYER MET2 ;
      RECT 4.9 4.75 5.4 5.15 ;
      RECT 3.35 4.75 3.75 5.15 ;
      RECT 3.3 4.8 5.4 5.1 ;
      RECT 3.3 2.85 3.8 3.25 ;
      RECT 1.35 2.85 1.85 3.25 ;
      RECT 1.35 2.9 3.8 3.2 ;
    LAYER VIA12 ;
      RECT 5.02 4.82 5.28 5.08 ;
      RECT 3.42 2.92 3.68 3.18 ;
      RECT 3.42 4.82 3.68 5.08 ;
      RECT 1.47 2.92 1.73 3.18 ;
    LAYER MET1 ;
      RECT 4.05 0.95 4.35 7.15 ;
      RECT 3.6 4 4.35 4.45 ;
      RECT 2.25 0.95 2.55 7.15 ;
      RECT 3.35 4.75 3.8 5.2 ;
      RECT 2.25 4.8 3.8 5.1 ;
      RECT 1.45 0.95 1.75 7.15 ;
      RECT 1.35 2.9 1.85 3.2 ;
      RECT 4.9 4.8 5.4 5.1 ;
      RECT 3.3 2.9 3.8 3.2 ;
  END
END gf180mcu_osu_sc_12T_lshifup
