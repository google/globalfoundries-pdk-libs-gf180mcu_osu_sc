# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_12T_dff_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN gf180mcu_osu_sc_12T_dff_1 0 -0.15 ;
  SIZE 13 BY 8.1 ;
  SYMMETRY X Y ;
  SITE GF018hv5v_mcu_sc7 ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER MET1 ;
        RECT 7.65 4 8.15 4.3 ;
        RECT 5.5 4 6.55 4.3 ;
        RECT 5.4 2 5.9 2.3 ;
        RECT 5.5 2 5.8 4.3 ;
        RECT 2.6 4 3.75 4.3 ;
        RECT 3.25 2.05 3.75 2.35 ;
        RECT 3.35 2.05 3.65 4.3 ;
      LAYER MET2 ;
        RECT 3.25 4 8.15 4.3 ;
        RECT 7.7 3.95 8.1 4.35 ;
        RECT 6.05 3.95 6.55 4.35 ;
        RECT 3.25 3.95 3.7 4.35 ;
      LAYER VIA12 ;
        RECT 3.37 4.02 3.63 4.28 ;
        RECT 6.17 4.02 6.43 4.28 ;
        RECT 7.77 4.02 8.03 4.28 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.9 3.35 2.4 3.65 ;
      LAYER MET2 ;
        RECT 1.75 3.35 2.55 3.65 ;
        RECT 1.9 3.3 2.4 3.7 ;
      LAYER VIA12 ;
        RECT 2.02 3.37 2.28 3.63 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 12.15 4.65 12.65 5 ;
        RECT 12.15 4.6 12.6 5 ;
        RECT 12.15 0.8 12.4 7 ;
      LAYER MET2 ;
        RECT 12.15 4.65 12.65 4.95 ;
        RECT 12.2 4.6 12.6 5 ;
      LAYER VIA12 ;
        RECT 12.27 4.67 12.53 4.93 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 10.45 4 11.9 4.3 ;
        RECT 11.55 1.9 11.8 4.3 ;
        RECT 10.45 1.9 11.8 2.15 ;
        RECT 10.45 4 10.7 7 ;
        RECT 10.45 0.8 10.7 2.15 ;
      LAYER MET2 ;
        RECT 11.4 4 11.9 4.3 ;
        RECT 11.45 3.95 11.85 4.35 ;
      LAYER VIA12 ;
        RECT 11.52 4.02 11.78 4.28 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.35 13 7.95 ;
        RECT 11.3 5.3 11.55 7.95 ;
        RECT 8.85 5.3 9.1 7.95 ;
        RECT 7.25 6.05 7.5 7.95 ;
        RECT 4.45 5.3 4.7 7.95 ;
        RECT 1.4 5.3 1.65 7.95 ;
      LAYER MET2 ;
        RECT 11.25 7.4 11.75 7.7 ;
        RECT 11.3 7.35 11.7 7.75 ;
        RECT 10.05 7.4 10.55 7.7 ;
        RECT 10.1 7.35 10.5 7.75 ;
        RECT 8.85 7.4 9.35 7.7 ;
        RECT 8.9 7.35 9.3 7.75 ;
        RECT 7.65 7.4 8.15 7.7 ;
        RECT 7.7 7.35 8.1 7.75 ;
        RECT 6.45 7.4 6.95 7.7 ;
        RECT 6.5 7.35 6.9 7.75 ;
        RECT 5.25 7.4 5.75 7.7 ;
        RECT 5.3 7.35 5.7 7.75 ;
        RECT 4.05 7.4 4.55 7.7 ;
        RECT 4.1 7.35 4.5 7.75 ;
        RECT 2.85 7.4 3.35 7.7 ;
        RECT 2.9 7.35 3.3 7.75 ;
        RECT 1.65 7.4 2.15 7.7 ;
        RECT 1.7 7.35 2.1 7.75 ;
        RECT 0.45 7.4 0.95 7.7 ;
        RECT 0.5 7.35 0.9 7.75 ;
      LAYER VIA12 ;
        RECT 0.57 7.42 0.83 7.68 ;
        RECT 1.77 7.42 2.03 7.68 ;
        RECT 2.97 7.42 3.23 7.68 ;
        RECT 4.17 7.42 4.43 7.68 ;
        RECT 5.37 7.42 5.63 7.68 ;
        RECT 6.57 7.42 6.83 7.68 ;
        RECT 7.77 7.42 8.03 7.68 ;
        RECT 8.97 7.42 9.23 7.68 ;
        RECT 10.17 7.42 10.43 7.68 ;
        RECT 11.37 7.42 11.63 7.68 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 -0.15 13 0.45 ;
        RECT 11.3 -0.15 11.55 1.65 ;
        RECT 8.85 -0.15 9.1 1.3 ;
        RECT 7.25 -0.15 7.5 1.65 ;
        RECT 4.45 -0.15 4.7 1.25 ;
        RECT 1.4 -0.15 1.65 1.65 ;
      LAYER MET2 ;
        RECT 11.25 0.1 11.75 0.4 ;
        RECT 11.3 0.05 11.7 0.45 ;
        RECT 10.05 0.1 10.55 0.4 ;
        RECT 10.1 0.05 10.5 0.45 ;
        RECT 8.85 0.1 9.35 0.4 ;
        RECT 8.9 0.05 9.3 0.45 ;
        RECT 7.65 0.1 8.15 0.4 ;
        RECT 7.7 0.05 8.1 0.45 ;
        RECT 6.45 0.1 6.95 0.4 ;
        RECT 6.5 0.05 6.9 0.45 ;
        RECT 5.25 0.1 5.75 0.4 ;
        RECT 5.3 0.05 5.7 0.45 ;
        RECT 4.05 0.1 4.55 0.4 ;
        RECT 4.1 0.05 4.5 0.45 ;
        RECT 2.85 0.1 3.35 0.4 ;
        RECT 2.9 0.05 3.3 0.45 ;
        RECT 1.65 0.1 2.15 0.4 ;
        RECT 1.7 0.05 2.1 0.45 ;
        RECT 0.45 0.1 0.95 0.4 ;
        RECT 0.5 0.05 0.9 0.45 ;
      LAYER VIA12 ;
        RECT 0.57 0.12 0.83 0.38 ;
        RECT 1.77 0.12 2.03 0.38 ;
        RECT 2.97 0.12 3.23 0.38 ;
        RECT 4.17 0.12 4.43 0.38 ;
        RECT 5.37 0.12 5.63 0.38 ;
        RECT 6.57 0.12 6.83 0.38 ;
        RECT 7.77 0.12 8.03 0.38 ;
        RECT 8.97 0.12 9.23 0.38 ;
        RECT 10.17 0.12 10.43 0.38 ;
        RECT 11.37 0.12 11.63 0.38 ;
    END
  END VSS
  OBS
    LAYER MET2 ;
      RECT 6.75 4.6 7.15 5 ;
      RECT 6.7 4.65 9.9 4.95 ;
      RECT 9.6 2.7 9.9 4.95 ;
      RECT 10.7 2.65 11.1 3.05 ;
      RECT 9.6 2.7 11.15 3 ;
      RECT 9 1.5 9.4 1.9 ;
      RECT 8.5 1.55 9.45 1.85 ;
      RECT 5.8 1.35 6.2 1.75 ;
      RECT 5.75 1.4 8.8 1.7 ;
      RECT 5.75 1.5 9.4 1.7 ;
      RECT 8.05 2.65 8.45 3.05 ;
      RECT 6.1 2.65 6.5 3.05 ;
      RECT 6.05 2.7 8.55 3 ;
      RECT 6.8 3.3 7.2 3.7 ;
      RECT 6.75 3.35 7.25 3.65 ;
      RECT 4.1 2 4.5 2.4 ;
      RECT 0.45 2 0.85 2.4 ;
      RECT 0.4 2.05 4.55 2.35 ;
    LAYER VIA12 ;
      RECT 10.77 2.72 11.03 2.98 ;
      RECT 9.07 1.57 9.33 1.83 ;
      RECT 8.12 2.72 8.38 2.98 ;
      RECT 6.87 3.37 7.13 3.63 ;
      RECT 6.82 4.67 7.08 4.93 ;
      RECT 6.17 2.72 6.43 2.98 ;
      RECT 5.87 1.42 6.13 1.68 ;
      RECT 4.17 2.07 4.43 2.33 ;
      RECT 0.52 2.07 0.78 2.33 ;
    LAYER MET1 ;
      RECT 9.7 0.8 9.95 7 ;
      RECT 9.7 2.7 11.15 3 ;
      RECT 9.05 1.55 9.35 3.1 ;
      RECT 8.95 2.7 9.45 3 ;
      RECT 8.95 1.55 9.45 1.85 ;
      RECT 8.1 4.6 8.35 7 ;
      RECT 8.1 4.6 8.9 4.85 ;
      RECT 8.6 3.4 8.9 4.85 ;
      RECT 8.1 3.4 8.9 3.65 ;
      RECT 8.1 2.6 8.4 3.65 ;
      RECT 8.1 0.8 8.35 3.65 ;
      RECT 6.7 4.65 7.2 4.95 ;
      RECT 6.8 3.3 7.1 4.95 ;
      RECT 6.75 3.35 7.3 3.65 ;
      RECT 6.8 3.3 7.2 3.65 ;
      RECT 5.85 5.8 6.1 7 ;
      RECT 4.95 5.8 6.1 6.05 ;
      RECT 4.95 3.3 5.2 6.05 ;
      RECT 4.9 1.45 5.15 3.55 ;
      RECT 4.9 1.45 6.25 1.7 ;
      RECT 5.85 1.4 6.25 1.7 ;
      RECT 5.85 0.8 6.1 1.7 ;
      RECT 4.05 4.65 4.55 4.95 ;
      RECT 4.15 2.05 4.45 4.95 ;
      RECT 4.05 2.05 4.55 2.35 ;
      RECT 3.05 4.8 3.3 7 ;
      RECT 1.4 4.8 3.3 5.05 ;
      RECT 1.4 2.1 1.65 5.05 ;
      RECT 1.05 4 1.65 4.3 ;
      RECT 1.4 2.1 2.4 2.35 ;
      RECT 2 1.4 2.4 2.35 ;
      RECT 2 1.4 3.3 1.65 ;
      RECT 3.05 0.8 3.3 1.65 ;
      RECT 0.55 0.8 0.8 7 ;
      RECT 0.5 1.95 0.8 2.45 ;
      RECT 6.05 2.7 6.55 3 ;
  END
END gf180mcu_osu_sc_12T_dff_1
