magic
tech gf180mcuC
timestamp 1661875423
<< nwell >>
rect 0 61 76 123
<< nmos >>
rect 16 19 22 36
rect 33 19 39 36
rect 50 19 56 36
<< pmos >>
rect 19 70 25 104
rect 30 70 36 104
rect 50 70 56 104
<< ndiff >>
rect 6 27 16 36
rect 6 21 8 27
rect 13 21 16 27
rect 6 19 16 21
rect 22 32 33 36
rect 22 21 25 32
rect 30 21 33 32
rect 22 19 33 21
rect 39 34 50 36
rect 39 21 42 34
rect 47 21 50 34
rect 39 19 50 21
rect 56 34 66 36
rect 56 21 59 34
rect 64 21 66 34
rect 56 19 66 21
<< pdiff >>
rect 9 102 19 104
rect 9 72 11 102
rect 16 72 19 102
rect 9 70 19 72
rect 25 70 30 104
rect 36 102 50 104
rect 36 88 39 102
rect 47 88 50 102
rect 36 70 50 88
rect 56 102 66 104
rect 56 88 59 102
rect 64 88 66 102
rect 56 70 66 88
<< ndiffc >>
rect 8 21 13 27
rect 25 21 30 32
rect 42 21 47 34
rect 59 21 64 34
<< pdiffc >>
rect 11 72 16 102
rect 39 88 47 102
rect 59 88 64 102
<< psubdiff >>
rect 9 10 18 12
rect 9 5 11 10
rect 16 5 18 10
rect 9 3 18 5
rect 33 10 42 12
rect 33 5 35 10
rect 40 5 42 10
rect 33 3 42 5
rect 57 10 66 12
rect 57 5 59 10
rect 64 5 66 10
rect 57 3 66 5
<< nsubdiff >>
rect 9 118 18 120
rect 9 113 11 118
rect 16 113 18 118
rect 9 111 18 113
rect 33 118 42 120
rect 33 113 35 118
rect 40 113 42 118
rect 33 111 42 113
rect 57 118 66 120
rect 57 113 59 118
rect 64 113 66 118
rect 57 111 66 113
<< psubdiffcont >>
rect 11 5 16 10
rect 35 5 40 10
rect 59 5 64 10
<< nsubdiffcont >>
rect 11 113 16 118
rect 35 113 40 118
rect 59 113 64 118
<< polysilicon >>
rect 19 104 25 109
rect 30 104 36 109
rect 50 104 56 109
rect 19 68 25 70
rect 16 63 25 68
rect 30 68 36 70
rect 30 65 39 68
rect 50 67 56 70
rect 49 65 59 67
rect 30 63 43 65
rect 16 52 22 63
rect 33 57 35 63
rect 41 57 43 63
rect 49 59 51 65
rect 57 59 59 65
rect 49 57 59 59
rect 33 55 43 57
rect 16 50 28 52
rect 16 44 20 50
rect 26 44 28 50
rect 16 42 28 44
rect 16 36 22 42
rect 33 36 39 55
rect 50 36 56 57
rect 16 14 22 19
rect 33 14 39 19
rect 50 14 56 19
<< polycontact >>
rect 35 57 41 63
rect 51 59 57 65
rect 20 44 26 50
<< metal1 >>
rect 0 118 76 123
rect 0 112 11 118
rect 17 112 35 118
rect 41 112 59 118
rect 65 112 76 118
rect 0 111 76 112
rect 11 102 16 104
rect 39 102 47 111
rect 39 86 47 88
rect 59 102 64 104
rect 16 75 54 81
rect 11 65 16 72
rect 8 59 16 65
rect 48 65 54 75
rect 59 76 64 88
rect 59 70 61 76
rect 67 70 69 76
rect 8 39 13 59
rect 33 57 35 63
rect 41 57 43 63
rect 48 59 51 65
rect 57 59 59 65
rect 18 44 20 50
rect 26 44 28 50
rect 8 34 30 39
rect 25 32 30 34
rect 8 27 13 29
rect 8 12 13 21
rect 25 19 30 21
rect 42 34 47 36
rect 42 12 47 21
rect 59 35 64 36
rect 59 34 61 35
rect 67 29 69 35
rect 59 19 64 21
rect 0 11 76 12
rect 0 5 11 11
rect 17 5 35 11
rect 41 5 59 11
rect 65 5 76 11
rect 0 0 76 5
<< via1 >>
rect 11 113 16 118
rect 16 113 17 118
rect 11 112 17 113
rect 35 113 40 118
rect 40 113 41 118
rect 35 112 41 113
rect 59 113 64 118
rect 64 113 65 118
rect 59 112 65 113
rect 61 70 67 76
rect 35 57 41 63
rect 20 44 26 50
rect 61 34 67 35
rect 61 29 64 34
rect 64 29 67 34
rect 11 10 17 11
rect 11 5 16 10
rect 16 5 17 10
rect 35 10 41 11
rect 35 5 40 10
rect 40 5 41 10
rect 59 10 65 11
rect 59 5 64 10
rect 64 5 65 10
<< metal2 >>
rect 9 118 19 119
rect 9 112 11 118
rect 17 112 19 118
rect 9 111 19 112
rect 33 118 43 119
rect 33 112 35 118
rect 41 112 43 118
rect 33 111 43 112
rect 57 118 67 119
rect 57 112 59 118
rect 65 112 67 118
rect 57 111 67 112
rect 59 76 69 77
rect 59 70 61 76
rect 67 70 69 76
rect 59 69 69 70
rect 33 63 43 64
rect 33 57 35 63
rect 41 57 43 63
rect 33 56 43 57
rect 18 50 28 51
rect 18 44 20 50
rect 26 44 28 50
rect 18 43 28 44
rect 61 36 67 69
rect 59 35 69 36
rect 59 29 61 35
rect 67 29 69 35
rect 59 28 69 29
rect 9 11 19 12
rect 9 5 11 11
rect 17 5 19 11
rect 9 4 19 5
rect 33 11 43 12
rect 33 5 35 11
rect 41 5 43 11
rect 33 4 43 5
rect 57 11 67 12
rect 57 5 59 11
rect 65 5 67 11
rect 57 4 67 5
<< labels >>
rlabel metal2 14 116 14 116 1 VDD
rlabel metal2 14 8 14 8 1 GND
rlabel metal2 23 47 23 47 1 A
port 2 n
rlabel metal2 38 60 38 60 1 B
port 1 n
rlabel metal2 64 73 64 73 1 Y
port 3 n
<< end >>
