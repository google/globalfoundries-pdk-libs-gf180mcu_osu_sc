# Copyright 2022 Google LLC
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#      http://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO gf180mcu_osu_sc_gp12t3v3__oai31_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN gf180mcu_osu_sc_gp12t3v3__oai31_1 0 0 ;
  SIZE 4.8 BY 8.1 ;
  SYMMETRY X Y ;
  SITE gf180mcu_osu_sc_gp12t3v3 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 7.5 4.8 8.1 ;
        RECT 3.85 5.45 4.1 8.1 ;
        RECT 1.05 5.45 1.3 8.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER MET1 ;
        RECT 0 0 4.8 0.6 ;
        RECT 2.25 0 2.5 1.5 ;
        RECT 0.55 0 0.8 1.8 ;
    END
  END VSS
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 0.95 2.85 1.45 3.15 ;
      LAYER MET2 ;
        RECT 0.95 2.8 1.45 3.2 ;
      LAYER VIA12 ;
        RECT 1.07 2.87 1.33 3.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 1.8 2.85 2.3 3.15 ;
      LAYER MET2 ;
        RECT 1.8 2.8 2.3 3.2 ;
      LAYER VIA12 ;
        RECT 1.92 2.87 2.18 3.13 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 2.55 4.15 3.05 4.45 ;
      LAYER MET2 ;
        RECT 2.55 4.1 3.05 4.5 ;
      LAYER VIA12 ;
        RECT 2.67 4.17 2.93 4.43 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3.1 2.85 3.6 3.15 ;
      LAYER MET2 ;
        RECT 3.1 2.8 3.6 3.2 ;
      LAYER VIA12 ;
        RECT 3.22 2.87 3.48 3.13 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER MET1 ;
        RECT 3 4.8 4.25 5.1 ;
        RECT 3.95 0.95 4.2 2.5 ;
        RECT 3.85 2.25 4.1 5.1 ;
        RECT 3 4.8 3.25 7.15 ;
      LAYER MET2 ;
        RECT 3.75 4.75 4.25 5.15 ;
      LAYER VIA12 ;
        RECT 3.87 4.82 4.13 5.08 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 1.4 1.75 3.35 2 ;
      RECT 3.1 0.95 3.35 2 ;
      RECT 1.4 0.95 1.65 2 ;
  END
END gf180mcu_osu_sc_gp12t3v3__oai31_1
